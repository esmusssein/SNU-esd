module xis (
	input		[7:0] data_in,
	output 	[31:0] data_out2
);
	reg [31:0] data_out = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
	
	assign data_out2 = data_out;
	
	always @ (*)begin
		case(data_in)
		0   : data_out <= 32'h0001d3bb; 1   : data_out <= 32'h0001b981; 2   : data_out <= 32'h0001a8fd; 3   : data_out <= 32'h00019cbe; 4   : data_out <= 32'h000192ee; 5   : data_out <= 32'h00018ab0; 6   : data_out <= 32'h00018390; 7   : data_out <= 32'h00017d42; 8   : data_out <= 32'h00017799; 9   : data_out <= 32'h00017272; 10  : data_out <= 32'h00016db6; 11  : data_out <= 32'h00016954; 12  : data_out <= 32'h0001653c; 13  : data_out <= 32'h00016166; 14  : data_out <= 32'h00015dc8; 15  : data_out <= 32'h00015a5c;
		16  : data_out <= 32'h0001571b; 17  : data_out <= 32'h00015401; 18  : data_out <= 32'h00015109; 19  : data_out <= 32'h00014e32; 20  : data_out <= 32'h00014b77; 21  : data_out <= 32'h000148d6; 22  : data_out <= 32'h0001464c; 23  : data_out <= 32'h000143d9; 24  : data_out <= 32'h0001417a; 25  : data_out <= 32'h00013f2d; 26  : data_out <= 32'h00013cf2; 27  : data_out <= 32'h00013ac7; 28  : data_out <= 32'h000138ab; 29  : data_out <= 32'h0001369d; 30  : data_out <= 32'h0001349c; 31  : data_out <= 32'h000132a7;
		32  : data_out <= 32'h000130be; 33  : data_out <= 32'h00012ee0; 34  : data_out <= 32'h00012d0d; 35  : data_out <= 32'h00012b43; 36  : data_out <= 32'h00012982; 37  : data_out <= 32'h000127cb; 38  : data_out <= 32'h0001261b; 39  : data_out <= 32'h00012474; 40  : data_out <= 32'h000122d4; 41  : data_out <= 32'h0001213b; 42  : data_out <= 32'h00011fa9; 43  : data_out <= 32'h00011e1e; 44  : data_out <= 32'h00011c99; 45  : data_out <= 32'h00011b1a; 46  : data_out <= 32'h000119a1; 47  : data_out <= 32'h0001182d;
		48  : data_out <= 32'h000116bf; 49  : data_out <= 32'h00011556; 50  : data_out <= 32'h000113f1; 51  : data_out <= 32'h00011292; 52  : data_out <= 32'h00011136; 53  : data_out <= 32'h00010fdf; 54  : data_out <= 32'h00010e8d; 55  : data_out <= 32'h00010d3e; 56  : data_out <= 32'h00010bf3; 57  : data_out <= 32'h00010aac; 58  : data_out <= 32'h00010969; 59  : data_out <= 32'h00010829; 60  : data_out <= 32'h000106ed; 61  : data_out <= 32'h000105b3; 62  : data_out <= 32'h0001047d; 63  : data_out <= 32'h0001034a;
		64  : data_out <= 32'h0001021a; 65  : data_out <= 32'h000100ed; 66  : data_out <= 32'h0000ffc2; 67  : data_out <= 32'h0000fe9b; 68  : data_out <= 32'h0000fd75; 69  : data_out <= 32'h0000fc53; 70  : data_out <= 32'h0000fb32; 71  : data_out <= 32'h0000fa15; 72  : data_out <= 32'h0000f8f9; 73  : data_out <= 32'h0000f7e0; 74  : data_out <= 32'h0000f6c9; 75  : data_out <= 32'h0000f5b4; 76  : data_out <= 32'h0000f4a1; 77  : data_out <= 32'h0000f390; 78  : data_out <= 32'h0000f280; 79  : data_out <= 32'h0000f173;
		80  : data_out <= 32'h0000f068; 81  : data_out <= 32'h0000ef5e; 82  : data_out <= 32'h0000ee56; 83  : data_out <= 32'h0000ed50; 84  : data_out <= 32'h0000ec4b; 85  : data_out <= 32'h0000eb48; 86  : data_out <= 32'h0000ea46; 87  : data_out <= 32'h0000e946; 88  : data_out <= 32'h0000e848; 89  : data_out <= 32'h0000e74a; 90  : data_out <= 32'h0000e64f; 91  : data_out <= 32'h0000e554; 92  : data_out <= 32'h0000e45b; 93  : data_out <= 32'h0000e363; 94  : data_out <= 32'h0000e26c; 95  : data_out <= 32'h0000e176;
		96  : data_out <= 32'h0000e082; 97  : data_out <= 32'h0000df8e; 98  : data_out <= 32'h0000de9c; 99  : data_out <= 32'h0000ddab; 100 : data_out <= 32'h0000dcbb; 101 : data_out <= 32'h0000dbcb; 102 : data_out <= 32'h0000dadd; 103 : data_out <= 32'h0000d9f0; 104 : data_out <= 32'h0000d903; 105 : data_out <= 32'h0000d818; 106 : data_out <= 32'h0000d72d; 107 : data_out <= 32'h0000d643; 108 : data_out <= 32'h0000d55a; 109 : data_out <= 32'h0000d472; 110 : data_out <= 32'h0000d38a; 111 : data_out <= 32'h0000d2a3;
		112 : data_out <= 32'h0000d1bd; 113 : data_out <= 32'h0000d0d8; 114 : data_out <= 32'h0000cff3; 115 : data_out <= 32'h0000cf0f; 116 : data_out <= 32'h0000ce2b; 117 : data_out <= 32'h0000cd48; 118 : data_out <= 32'h0000cc66; 119 : data_out <= 32'h0000cb84; 120 : data_out <= 32'h0000caa3; 121 : data_out <= 32'h0000c9c2; 122 : data_out <= 32'h0000c8e1; 123 : data_out <= 32'h0000c801; 124 : data_out <= 32'h0000c722; 125 : data_out <= 32'h0000c643; 126 : data_out <= 32'h0000c564; 127 : data_out <= 32'h0000c486;
		128 : data_out <= 32'h0000c3a8; 129 : data_out <= 32'h0000c2ca; 130 : data_out <= 32'h0000c1ed; 131 : data_out <= 32'h0000c110; 132 : data_out <= 32'h0000c033; 133 : data_out <= 32'h0000bf56; 134 : data_out <= 32'h0000be7a; 135 : data_out <= 32'h0000bd9e; 136 : data_out <= 32'h0000bcc2; 137 : data_out <= 32'h0000bbe6; 138 : data_out <= 32'h0000bb0b; 139 : data_out <= 32'h0000ba2f; 140 : data_out <= 32'h0000b954; 141 : data_out <= 32'h0000b879; 142 : data_out <= 32'h0000b79e; 143 : data_out <= 32'h0000b6c3;
		144 : data_out <= 32'h0000b5e8; 145 : data_out <= 32'h0000b50d; 146 : data_out <= 32'h0000b432; 147 : data_out <= 32'h0000b357; 148 : data_out <= 32'h0000b27c; 149 : data_out <= 32'h0000b1a0; 150 : data_out <= 32'h0000b0c5; 151 : data_out <= 32'h0000afea; 152 : data_out <= 32'h0000af0f; 153 : data_out <= 32'h0000ae33; 154 : data_out <= 32'h0000ad57; 155 : data_out <= 32'h0000ac7c; 156 : data_out <= 32'h0000aba0; 157 : data_out <= 32'h0000aac3; 158 : data_out <= 32'h0000a9e7; 159 : data_out <= 32'h0000a90a;
		160 : data_out <= 32'h0000a82d; 161 : data_out <= 32'h0000a750; 162 : data_out <= 32'h0000a672; 163 : data_out <= 32'h0000a594; 164 : data_out <= 32'h0000a4b5; 165 : data_out <= 32'h0000a3d6; 166 : data_out <= 32'h0000a2f7; 167 : data_out <= 32'h0000a218; 168 : data_out <= 32'h0000a137; 169 : data_out <= 32'h0000a057; 170 : data_out <= 32'h00009f75; 171 : data_out <= 32'h00009e94; 172 : data_out <= 32'h00009db1; 173 : data_out <= 32'h00009cce; 174 : data_out <= 32'h00009beb; 175 : data_out <= 32'h00009b07;
		176 : data_out <= 32'h00009a22; 177 : data_out <= 32'h0000993c; 178 : data_out <= 32'h00009856; 179 : data_out <= 32'h0000976e; 180 : data_out <= 32'h00009686; 181 : data_out <= 32'h0000959d; 182 : data_out <= 32'h000094b4; 183 : data_out <= 32'h000093c9; 184 : data_out <= 32'h000092dd; 185 : data_out <= 32'h000091f0; 186 : data_out <= 32'h00009103; 187 : data_out <= 32'h00009014; 188 : data_out <= 32'h00008f24; 189 : data_out <= 32'h00008e33; 190 : data_out <= 32'h00008d40; 191 : data_out <= 32'h00008c4d;
		192 : data_out <= 32'h00008b58; 193 : data_out <= 32'h00008a61; 194 : data_out <= 32'h0000896a; 195 : data_out <= 32'h00008871; 196 : data_out <= 32'h00008776; 197 : data_out <= 32'h00008679; 198 : data_out <= 32'h0000857b; 199 : data_out <= 32'h0000847c; 200 : data_out <= 32'h0000837a; 201 : data_out <= 32'h00008277; 202 : data_out <= 32'h00008172; 203 : data_out <= 32'h0000806a; 204 : data_out <= 32'h00007f61; 205 : data_out <= 32'h00007e55; 206 : data_out <= 32'h00007d47; 207 : data_out <= 32'h00007c37;
		208 : data_out <= 32'h00007b24; 209 : data_out <= 32'h00007a0f; 210 : data_out <= 32'h000078f7; 211 : data_out <= 32'h000077dc; 212 : data_out <= 32'h000076bf; 213 : data_out <= 32'h0000759e; 214 : data_out <= 32'h0000747a; 215 : data_out <= 32'h00007353; 216 : data_out <= 32'h00007228; 217 : data_out <= 32'h000070f9; 218 : data_out <= 32'h00006fc7; 219 : data_out <= 32'h00006e90; 220 : data_out <= 32'h00006d56; 221 : data_out <= 32'h00006c16; 222 : data_out <= 32'h00006ad2; 223 : data_out <= 32'h00006989;
		224 : data_out <= 32'h0000683b; 225 : data_out <= 32'h000066e7; 226 : data_out <= 32'h0000658d; 227 : data_out <= 32'h0000642c; 228 : data_out <= 32'h000062c5; 229 : data_out <= 32'h00006157; 230 : data_out <= 32'h00005fe1; 231 : data_out <= 32'h00005e62; 232 : data_out <= 32'h00005cdb; 233 : data_out <= 32'h00005b4a; 234 : data_out <= 32'h000059af; 235 : data_out <= 32'h00005808; 236 : data_out <= 32'h00005656; 237 : data_out <= 32'h00005495; 238 : data_out <= 32'h000052c6; 239 : data_out <= 32'h000050e7;
		240 : data_out <= 32'h00004ef6; 241 : data_out <= 32'h00004cf0; 242 : data_out <= 32'h00004ad4; 243 : data_out <= 32'h0000489e; 244 : data_out <= 32'h0000464a; 245 : data_out <= 32'h000043d4; 246 : data_out <= 32'h00004134; 247 : data_out <= 32'h00003e64; 248 : data_out <= 32'h00003b58; 249 : data_out <= 32'h00003800; 250 : data_out <= 32'h00003446; 251 : data_out <= 32'h00003003; 252 : data_out <= 32'h00002af9; 253 : data_out <= 32'h000024a1; 254 : data_out <= 32'h00001b8d; 255 : data_out <= 32'h00000000;			default: data_out <= 0;

		endcase
	end
endmodule

module yis (
	input		[7:0] data_in,
	output 	[31:0] data_out2
);
	reg [31:0] data_out = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
	
	assign data_out2 = data_out;
	
	always@(*)begin
		case(data_in)
		0   : data_out <= 32'h00000029; 1   : data_out <= 32'h00000055; 2   : data_out <= 32'h00000084; 3   : data_out <= 32'h000000b4; 4   : data_out <= 32'h000000e7; 5   : data_out <= 32'h0000011a; 6   : data_out <= 32'h0000014e; 7   : data_out <= 32'h00000184; 8   : data_out <= 32'h000001ba; 9   : data_out <= 32'h000001f1; 10  : data_out <= 32'h00000229; 11  : data_out <= 32'h00000261; 12  : data_out <= 32'h0000029a; 13  : data_out <= 32'h000002d4; 14  : data_out <= 32'h0000030f; 15  : data_out <= 32'h0000034a;
		16  : data_out <= 32'h00000386; 17  : data_out <= 32'h000003c2; 18  : data_out <= 32'h000003ff; 19  : data_out <= 32'h0000043c; 20  : data_out <= 32'h0000047a; 21  : data_out <= 32'h000004b8; 22  : data_out <= 32'h000004f7; 23  : data_out <= 32'h00000536; 24  : data_out <= 32'h00000576; 25  : data_out <= 32'h000005b6; 26  : data_out <= 32'h000005f7; 27  : data_out <= 32'h00000638; 28  : data_out <= 32'h0000067a; 29  : data_out <= 32'h000006bc; 30  : data_out <= 32'h000006ff; 31  : data_out <= 32'h00000742;
		32  : data_out <= 32'h00000785; 33  : data_out <= 32'h000007c9; 34  : data_out <= 32'h0000080d; 35  : data_out <= 32'h00000852; 36  : data_out <= 32'h00000897; 37  : data_out <= 32'h000008dd; 38  : data_out <= 32'h00000922; 39  : data_out <= 32'h00000969; 40  : data_out <= 32'h000009af; 41  : data_out <= 32'h000009f6; 42  : data_out <= 32'h00000a3e; 43  : data_out <= 32'h00000a86; 44  : data_out <= 32'h00000ace; 45  : data_out <= 32'h00000b17; 46  : data_out <= 32'h00000b60; 47  : data_out <= 32'h00000ba9;
		48  : data_out <= 32'h00000bf3; 49  : data_out <= 32'h00000c3d; 50  : data_out <= 32'h00000c88; 51  : data_out <= 32'h00000cd3; 52  : data_out <= 32'h00000d1e; 53  : data_out <= 32'h00000d69; 54  : data_out <= 32'h00000db5; 55  : data_out <= 32'h00000e02; 56  : data_out <= 32'h00000e4f; 57  : data_out <= 32'h00000e9c; 58  : data_out <= 32'h00000ee9; 59  : data_out <= 32'h00000f37; 60  : data_out <= 32'h00000f85; 61  : data_out <= 32'h00000fd4; 62  : data_out <= 32'h00001023; 63  : data_out <= 32'h00001072;
		64  : data_out <= 32'h000010c2; 65  : data_out <= 32'h00001112; 66  : data_out <= 32'h00001163; 67  : data_out <= 32'h000011b4; 68  : data_out <= 32'h00001205; 69  : data_out <= 32'h00001256; 70  : data_out <= 32'h000012a8; 71  : data_out <= 32'h000012fb; 72  : data_out <= 32'h0000134d; 73  : data_out <= 32'h000013a0; 74  : data_out <= 32'h000013f4; 75  : data_out <= 32'h00001447; 76  : data_out <= 32'h0000149c; 77  : data_out <= 32'h000014f0; 78  : data_out <= 32'h00001545; 79  : data_out <= 32'h0000159a;
		80  : data_out <= 32'h000015f0; 81  : data_out <= 32'h00001646; 82  : data_out <= 32'h0000169c; 83  : data_out <= 32'h000016f3; 84  : data_out <= 32'h0000174a; 85  : data_out <= 32'h000017a1; 86  : data_out <= 32'h000017f9; 87  : data_out <= 32'h00001852; 88  : data_out <= 32'h000018aa; 89  : data_out <= 32'h00001903; 90  : data_out <= 32'h0000195d; 91  : data_out <= 32'h000019b6; 92  : data_out <= 32'h00001a10; 93  : data_out <= 32'h00001a6b; 94  : data_out <= 32'h00001ac6; 95  : data_out <= 32'h00001b21;
		96  : data_out <= 32'h00001b7d; 97  : data_out <= 32'h00001bd9; 98  : data_out <= 32'h00001c35; 99  : data_out <= 32'h00001c92; 100 : data_out <= 32'h00001cf0; 101 : data_out <= 32'h00001d4d; 102 : data_out <= 32'h00001dab; 103 : data_out <= 32'h00001e0a; 104 : data_out <= 32'h00001e69; 105 : data_out <= 32'h00001ec8; 106 : data_out <= 32'h00001f27; 107 : data_out <= 32'h00001f88; 108 : data_out <= 32'h00001fe8; 109 : data_out <= 32'h00002049; 110 : data_out <= 32'h000020aa; 111 : data_out <= 32'h0000210c;
		112 : data_out <= 32'h0000216e; 113 : data_out <= 32'h000021d1; 114 : data_out <= 32'h00002234; 115 : data_out <= 32'h00002297; 116 : data_out <= 32'h000022fb; 117 : data_out <= 32'h0000235f; 118 : data_out <= 32'h000023c4; 119 : data_out <= 32'h00002429; 120 : data_out <= 32'h0000248f; 121 : data_out <= 32'h000024f5; 122 : data_out <= 32'h0000255b; 123 : data_out <= 32'h000025c2; 124 : data_out <= 32'h00002629; 125 : data_out <= 32'h00002691; 126 : data_out <= 32'h000026f9; 127 : data_out <= 32'h00002762;
		128 : data_out <= 32'h000027cb; 129 : data_out <= 32'h00002835; 130 : data_out <= 32'h0000289f; 131 : data_out <= 32'h0000290a; 132 : data_out <= 32'h00002975; 133 : data_out <= 32'h000029e0; 134 : data_out <= 32'h00002a4c; 135 : data_out <= 32'h00002ab9; 136 : data_out <= 32'h00002b26; 137 : data_out <= 32'h00002b93; 138 : data_out <= 32'h00002c01; 139 : data_out <= 32'h00002c70; 140 : data_out <= 32'h00002cdf; 141 : data_out <= 32'h00002d4f; 142 : data_out <= 32'h00002dbf; 143 : data_out <= 32'h00002e2f;
		144 : data_out <= 32'h00002ea0; 145 : data_out <= 32'h00002f12; 146 : data_out <= 32'h00002f84; 147 : data_out <= 32'h00002ff7; 148 : data_out <= 32'h0000306a; 149 : data_out <= 32'h000030de; 150 : data_out <= 32'h00003152; 151 : data_out <= 32'h000031c7; 152 : data_out <= 32'h0000323d; 153 : data_out <= 32'h000032b3; 154 : data_out <= 32'h0000332a; 155 : data_out <= 32'h000033a1; 156 : data_out <= 32'h00003419; 157 : data_out <= 32'h00003491; 158 : data_out <= 32'h0000350a; 159 : data_out <= 32'h00003584;
		160 : data_out <= 32'h000035fe; 161 : data_out <= 32'h00003679; 162 : data_out <= 32'h000036f5; 163 : data_out <= 32'h00003771; 164 : data_out <= 32'h000037ee; 165 : data_out <= 32'h0000386b; 166 : data_out <= 32'h000038e9; 167 : data_out <= 32'h00003968; 168 : data_out <= 32'h000039e8; 169 : data_out <= 32'h00003a68; 170 : data_out <= 32'h00003ae9; 171 : data_out <= 32'h00003b6a; 172 : data_out <= 32'h00003bed; 173 : data_out <= 32'h00003c70; 174 : data_out <= 32'h00003cf4; 175 : data_out <= 32'h00003d78;
		176 : data_out <= 32'h00003dfe; 177 : data_out <= 32'h00003e84; 178 : data_out <= 32'h00003f0b; 179 : data_out <= 32'h00003f92; 180 : data_out <= 32'h0000401b; 181 : data_out <= 32'h000040a4; 182 : data_out <= 32'h0000412e; 183 : data_out <= 32'h000041b9; 184 : data_out <= 32'h00004245; 185 : data_out <= 32'h000042d2; 186 : data_out <= 32'h00004360; 187 : data_out <= 32'h000043ee; 188 : data_out <= 32'h0000447e; 189 : data_out <= 32'h0000450e; 190 : data_out <= 32'h000045a0; 191 : data_out <= 32'h00004632;
		192 : data_out <= 32'h000046c5; 193 : data_out <= 32'h0000475a; 194 : data_out <= 32'h000047ef; 195 : data_out <= 32'h00004885; 196 : data_out <= 32'h0000491d; 197 : data_out <= 32'h000049b6; 198 : data_out <= 32'h00004a4f; 199 : data_out <= 32'h00004aea; 200 : data_out <= 32'h00004b86; 201 : data_out <= 32'h00004c23; 202 : data_out <= 32'h00004cc2; 203 : data_out <= 32'h00004d62; 204 : data_out <= 32'h00004e03; 205 : data_out <= 32'h00004ea5; 206 : data_out <= 32'h00004f48; 207 : data_out <= 32'h00004fed;
		208 : data_out <= 32'h00005094; 209 : data_out <= 32'h0000513c; 210 : data_out <= 32'h000051e5; 211 : data_out <= 32'h00005290; 212 : data_out <= 32'h0000533c; 213 : data_out <= 32'h000053eb; 214 : data_out <= 32'h0000549a; 215 : data_out <= 32'h0000554c; 216 : data_out <= 32'h000055ff; 217 : data_out <= 32'h000056b4; 218 : data_out <= 32'h0000576b; 219 : data_out <= 32'h00005824; 220 : data_out <= 32'h000058df; 221 : data_out <= 32'h0000599c; 222 : data_out <= 32'h00005a5b; 223 : data_out <= 32'h00005b1d;
		224 : data_out <= 32'h00005be1; 225 : data_out <= 32'h00005ca7; 226 : data_out <= 32'h00005d70; 227 : data_out <= 32'h00005e3c; 228 : data_out <= 32'h00005f0a; 229 : data_out <= 32'h00005fdb; 230 : data_out <= 32'h000060b0; 231 : data_out <= 32'h00006187; 232 : data_out <= 32'h00006262; 233 : data_out <= 32'h00006341; 234 : data_out <= 32'h00006423; 235 : data_out <= 32'h0000650a; 236 : data_out <= 32'h000065f5; 237 : data_out <= 32'h000066e4; 238 : data_out <= 32'h000067d8; 239 : data_out <= 32'h000068d2;
		240 : data_out <= 32'h000069d2; 241 : data_out <= 32'h00006ad7; 242 : data_out <= 32'h00006be4; 243 : data_out <= 32'h00006cf8; 244 : data_out <= 32'h00006e15; 245 : data_out <= 32'h00006f3b; 246 : data_out <= 32'h0000706c; 247 : data_out <= 32'h000071a9; 248 : data_out <= 32'h000072f4; 249 : data_out <= 32'h00007451; 250 : data_out <= 32'h000075c2; 251 : data_out <= 32'h0000774d; 252 : data_out <= 32'h000078fc; 253 : data_out <= 32'h00007add; 254 : data_out <= 32'h00007d11; 255 : data_out <= 32'h00008000;
		endcase
	end
endmodule


module sqrt_minus2_ln (
	input		[14:0] data_in;
	output 	[31:0] data_out;
);
	always@(*)begin
		case(data_in)
		default:
		endcase
	end
endmodule

module cosin (
	input		[14:0] data_in;
	output 	[31:0] data_out;
);
	always@(*)begin
		case(data_in)
		default:
		endcase
	end
endmodule

module sin (
	input		[14:0] data_in;
	output 	[31:0] data_out;
);
	always@(*)begin
		case(data_in)
		default:
		endcase
	end
endmodule
		
// megafunction wizard: %RAM initializer%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTMEM_INIT 

// ============================================================
// File Name: ram.v
// Megafunction Name(s):
// 			ALTMEM_INIT
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 11.0 Build 157 04/27/2011 SJ Web Edition
// ************************************************************

//Copyright (C) 1991-2011 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.

module ram (
	clock,
	init,
	dataout,
	init_busy,
	ram_address,
	ram_wren)/* synthesis synthesis_clearbox = 1 */;

	input	  clock;
	input	  init;
	output	[31:0]  dataout;
	output	  init_busy;
	output	[16:0]  ram_address;
	output	  ram_wren;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
// Retrieval info: CONSTANT: INIT_FILE STRING "UNUSED"
// Retrieval info: CONSTANT: INIT_TO_ZERO STRING "YES"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
// Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altmem_init"
// Retrieval info: CONSTANT: NUMWORDS NUMERIC "100000"
// Retrieval info: CONSTANT: PORT_ROM_DATA_READY STRING "PORT_UNUSED"
// Retrieval info: CONSTANT: ROM_READ_LATENCY NUMERIC "1"
// Retrieval info: CONSTANT: WIDTH NUMERIC "32"
// Retrieval info: CONSTANT: WIDTHAD NUMERIC "17"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: USED_PORT: dataout 0 0 32 0 OUTPUT NODEFVAL "dataout[31..0]"
// Retrieval info: CONNECT: dataout 0 0 32 0 @dataout 0 0 32 0
// Retrieval info: USED_PORT: init 0 0 0 0 INPUT NODEFVAL "init"
// Retrieval info: CONNECT: @init 0 0 0 0 init 0 0 0 0
// Retrieval info: USED_PORT: init_busy 0 0 0 0 OUTPUT NODEFVAL "init_busy"
// Retrieval info: CONNECT: init_busy 0 0 0 0 @init_busy 0 0 0 0
// Retrieval info: USED_PORT: ram_address 0 0 17 0 OUTPUT NODEFVAL "ram_address[16..0]"
// Retrieval info: CONNECT: ram_address 0 0 17 0 @ram_address 0 0 17 0
// Retrieval info: USED_PORT: ram_wren 0 0 0 0 OUTPUT NODEFVAL "ram_wren"
// Retrieval info: CONNECT: ram_wren 0 0 0 0 @ram_wren 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL ram.v TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL ram.qip TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL ram.bsf TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ram_inst.v TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ram_bb.v TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ram.inc TRUE TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL ram.cmp TRUE TRUE
// Retrieval info: LIB_FILE: lpm

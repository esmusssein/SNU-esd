module cosin (
	input	[7:0] data_in,
	output [14:0] cos_x_out
);

	reg [31:0] x = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
	
	assign cos_x_out = x;
	
	always @(*) begin
		case(data_in)
		10'h  1: x = 16'hffff; 10'h  2: x = 16'hfffe; 10'h  3: x = 16'hfffd; 10'h  4: x = 16'hfffb; 10'h  5: x = 16'hfff8; 10'h  6: x = 16'hfff4; 10'h  7: x = 16'hfff0; 10'h  8: x = 16'hffec; 10'h  9: x = 16'hffe7; 10'h  a: x = 16'hffe1; 10'h  b: x = 16'hffda; 10'h  c: x = 16'hffd3; 10'h  d: x = 16'hffcb; 10'h  e: x = 16'hffc3; 10'h  f: x = 16'hffba; 10'h 10: x = 16'hffb1; 10'h 11: x = 16'hffa6; 10'h 12: x = 16'hff9c; 10'h 13: x = 16'hff90; 10'h 14: x = 16'hff84; 10'h 15: x = 16'hff78; 10'h 16: x = 16'hff6a; 10'h 17: x = 16'hff5c; 10'h 18: x = 16'hff4e; 10'h 19: x = 16'hff3f; 10'h 1a: x = 16'hff2f; 10'h 1b: x = 16'hff1f; 10'h 1c: x = 16'hff0e; 10'h 1d: x = 16'hfefc; 10'h 1e: x = 16'hfeea; 10'h 1f: x = 16'hfed7; 10'h 20: x = 16'hfec4; 10'h 21: x = 16'hfeb0; 10'h 22: x = 16'hfe9b; 10'h 23: x = 16'hfe86; 10'h 24: x = 16'hfe70; 10'h 25: x = 16'hfe5a; 10'h 26: x = 16'hfe43; 10'h 27: x = 16'hfe2b; 10'h 28: x = 16'hfe13; 10'h 29: x = 16'hfdfa; 10'h 2a: x = 16'hfde0; 10'h 2b: x = 16'hfdc6; 10'h 2c: x = 16'hfdab; 10'h 2d: x = 16'hfd90; 10'h 2e: x = 16'hfd74; 10'h 2f: x = 16'hfd57; 10'h 30: x = 16'hfd3a; 10'h 31: x = 16'hfd1c; 10'h 32: x = 16'hfcfe; 10'h 33: x = 16'hfcdf; 10'h 34: x = 16'hfcbf; 10'h 35: x = 16'hfc9f; 10'h 36: x = 16'hfc7e; 10'h 37: x = 16'hfc5d; 10'h 38: x = 16'hfc3b; 10'h 39: x = 16'hfc18; 10'h 3a: x = 16'hfbf5; 10'h 3b: x = 16'hfbd1; 10'h 3c: x = 16'hfbac; 10'h 3d: x = 16'hfb87; 10'h 3e: x = 16'hfb61; 10'h 3f: x = 16'hfb3b; 10'h 40: x = 16'hfb14; 10'h 41: x = 16'hfaed; 10'h 42: x = 16'hfac5; 10'h 43: x = 16'hfa9c; 10'h 44: x = 16'hfa73; 10'h 45: x = 16'hfa49; 10'h 46: x = 16'hfa1e; 10'h 47: x = 16'hf9f3; 10'h 48: x = 16'hf9c7; 10'h 49: x = 16'hf99b; 10'h 4a: x = 16'hf96e; 10'h 4b: x = 16'hf940; 10'h 4c: x = 16'hf912; 10'h 4d: x = 16'hf8e3; 10'h 4e: x = 16'hf8b4; 10'h 4f: x = 16'hf884; 10'h 50: x = 16'hf853; 10'h 51: x = 16'hf822; 10'h 52: x = 16'hf7f1; 10'h 53: x = 16'hf7be; 10'h 54: x = 16'hf78b; 10'h 55: x = 16'hf758; 10'h 56: x = 16'hf724; 10'h 57: x = 16'hf6ef; 10'h 58: x = 16'hf6ba; 10'h 59: x = 16'hf684; 10'h 5a: x = 16'hf64d; 10'h 5b: x = 16'hf616; 10'h 5c: x = 16'hf5de; 10'h 5d: x = 16'hf5a6; 10'h 5e: x = 16'hf56d; 10'h 5f: x = 16'hf534; 10'h 60: x = 16'hf4fa; 10'h 61: x = 16'hf4bf; 10'h 62: x = 16'hf484; 10'h 63: x = 16'hf448; 10'h 64: x = 16'hf40b; 10'h 65: x = 16'hf3ce; 10'h 66: x = 16'hf391; 10'h 67: x = 16'hf353; 10'h 68: x = 16'hf314; 10'h 69: x = 16'hf2d4; 10'h 6a: x = 16'hf294; 10'h 6b: x = 16'hf254; 10'h 6c: x = 16'hf213; 10'h 6d: x = 16'hf1d1; 10'h 6e: x = 16'hf18f; 10'h 6f: x = 16'hf14c; 10'h 70: x = 16'hf109; 10'h 71: x = 16'hf0c5; 10'h 72: x = 16'hf080; 10'h 73: x = 16'hf03b; 10'h 74: x = 16'heff5; 10'h 75: x = 16'hefaf; 10'h 76: x = 16'hef68; 10'h 77: x = 16'hef20; 10'h 78: x = 16'heed8; 10'h 79: x = 16'hee8f; 10'h 7a: x = 16'hee46; 10'h 7b: x = 16'hedfc; 10'h 7c: x = 16'hedb2; 10'h 7d: x = 16'hed67; 10'h 7e: x = 16'hed1c; 10'h 7f: x = 16'hecd0; 10'h 80: x = 16'hec83; 10'h 81: x = 16'hec36; 10'h 82: x = 16'hebe8; 10'h 83: x = 16'heb99; 10'h 84: x = 16'heb4b; 10'h 85: x = 16'heafb; 10'h 86: x = 16'heaab; 10'h 87: x = 16'hea5a; 10'h 88: x = 16'hea09; 10'h 89: x = 16'he9b7; 10'h 8a: x = 16'he965; 10'h 8b: x = 16'he912; 10'h 8c: x = 16'he8bf; 10'h 8d: x = 16'he86b; 10'h 8e: x = 16'he816; 10'h 8f: x = 16'he7c1; 10'h 90: x = 16'he76b; 10'h 91: x = 16'he715; 10'h 92: x = 16'he6be; 10'h 93: x = 16'he667; 10'h 94: x = 16'he60f; 10'h 95: x = 16'he5b7; 10'h 96: x = 16'he55e; 10'h 97: x = 16'he504; 10'h 98: x = 16'he4aa; 10'h 99: x = 16'he44f; 10'h 9a: x = 16'he3f4; 10'h 9b: x = 16'he398; 10'h 9c: x = 16'he33c; 10'h 9d: x = 16'he2df; 10'h 9e: x = 16'he282; 10'h 9f: x = 16'he224; 10'h a0: x = 16'he1c5; 10'h a1: x = 16'he166; 10'h a2: x = 16'he106; 10'h a3: x = 16'he0a6; 10'h a4: x = 16'he046; 10'h a5: x = 16'hdfe4; 10'h a6: x = 16'hdf83; 10'h a7: x = 16'hdf20; 10'h a8: x = 16'hdebe; 10'h a9: x = 16'hde5a; 10'h aa: x = 16'hddf6; 10'h ab: x = 16'hdd92; 10'h ac: x = 16'hdd2d; 10'h ad: x = 16'hdcc7; 10'h ae: x = 16'hdc61; 10'h af: x = 16'hdbfb; 10'h b0: x = 16'hdb94; 10'h b1: x = 16'hdb2c; 10'h b2: x = 16'hdac4; 10'h b3: x = 16'hda5b; 10'h b4: x = 16'hd9f2; 10'h b5: x = 16'hd988; 10'h b6: x = 16'hd91e; 10'h b7: x = 16'hd8b3; 10'h b8: x = 16'hd848; 10'h b9: x = 16'hd7dc; 10'h ba: x = 16'hd770; 10'h bb: x = 16'hd703; 10'h bc: x = 16'hd695; 10'h bd: x = 16'hd627; 10'h be: x = 16'hd5b9; 10'h bf: x = 16'hd54a; 10'h c0: x = 16'hd4db; 10'h c1: x = 16'hd46b; 10'h c2: x = 16'hd3fa; 10'h c3: x = 16'hd389; 10'h c4: x = 16'hd318; 10'h c5: x = 16'hd2a6; 10'h c6: x = 16'hd233; 10'h c7: x = 16'hd1c0; 10'h c8: x = 16'hd14d; 10'h c9: x = 16'hd0d9; 10'h ca: x = 16'hd064; 10'h cb: x = 16'hcfef; 10'h cc: x = 16'hcf7a; 10'h cd: x = 16'hcf04; 10'h ce: x = 16'hce8d; 10'h cf: x = 16'hce16; 10'h d0: x = 16'hcd9f; 10'h d1: x = 16'hcd26; 10'h d2: x = 16'hccae; 10'h d3: x = 16'hcc35; 10'h d4: x = 16'hcbbb; 10'h d5: x = 16'hcb41; 10'h d6: x = 16'hcac7; 10'h d7: x = 16'hca4c; 10'h d8: x = 16'hc9d1; 10'h d9: x = 16'hc955; 10'h da: x = 16'hc8d8; 10'h db: x = 16'hc85b; 10'h dc: x = 16'hc7de; 10'h dd: x = 16'hc760; 10'h de: x = 16'hc6e2; 10'h df: x = 16'hc663; 10'h e0: x = 16'hc5e4; 10'h e1: x = 16'hc564; 10'h e2: x = 16'hc4e3; 10'h e3: x = 16'hc463; 10'h e4: x = 16'hc3e2; 10'h e5: x = 16'hc360; 10'h e6: x = 16'hc2de; 10'h e7: x = 16'hc25b; 10'h e8: x = 16'hc1d8; 10'h e9: x = 16'hc154; 10'h ea: x = 16'hc0d0; 10'h eb: x = 16'hc04c; 10'h ec: x = 16'hbfc7; 10'h ed: x = 16'hbf41; 10'h ee: x = 16'hbebc; 10'h ef: x = 16'hbe35; 10'h f0: x = 16'hbdae; 10'h f1: x = 16'hbd27; 10'h f2: x = 16'hbca0; 10'h f3: x = 16'hbc17; 10'h f4: x = 16'hbb8f; 10'h f5: x = 16'hbb06; 10'h f6: x = 16'hba7c; 10'h f7: x = 16'hb9f2; 10'h f8: x = 16'hb968; 10'h f9: x = 16'hb8dd; 10'h fa: x = 16'hb852; 10'h fb: x = 16'hb7c6; 10'h fc: x = 16'hb73a; 10'h fd: x = 16'hb6ad; 10'h fe: x = 16'hb620; 10'h ff: x = 16'hb592; 10'h100: x = 16'hb504; 10'h101: x = 16'hb476; 10'h102: x = 16'hb3e7; 10'h103: x = 16'hb358; 10'h104: x = 16'hb2c8; 10'h105: x = 16'hb238; 10'h106: x = 16'hb1a8; 10'h107: x = 16'hb117; 10'h108: x = 16'hb085; 10'h109: x = 16'haff3; 10'h10a: x = 16'haf61; 10'h10b: x = 16'haece; 10'h10c: x = 16'hae3b; 10'h10d: x = 16'hada8; 10'h10e: x = 16'had14; 10'h10f: x = 16'hac80; 10'h110: x = 16'habeb; 10'h111: x = 16'hab56; 10'h112: x = 16'haac0; 10'h113: x = 16'haa2a; 10'h114: x = 16'ha994; 10'h115: x = 16'ha8fd; 10'h116: x = 16'ha866; 10'h117: x = 16'ha7ce; 10'h118: x = 16'ha736; 10'h119: x = 16'ha69d; 10'h11a: x = 16'ha605; 10'h11b: x = 16'ha56b; 10'h11c: x = 16'ha4d2; 10'h11d: x = 16'ha438; 10'h11e: x = 16'ha39d; 10'h11f: x = 16'ha302; 10'h120: x = 16'ha267; 10'h121: x = 16'ha1cb; 10'h122: x = 16'ha12f; 10'h123: x = 16'ha093; 10'h124: x = 16'h9ff6; 10'h125: x = 16'h9f59; 10'h126: x = 16'h9ebc; 10'h127: x = 16'h9e1e; 10'h128: x = 16'h9d7f; 10'h129: x = 16'h9ce1; 10'h12a: x = 16'h9c42; 10'h12b: x = 16'h9ba2; 10'h12c: x = 16'h9b02; 10'h12d: x = 16'h9a62; 10'h12e: x = 16'h99c2; 10'h12f: x = 16'h9921; 10'h130: x = 16'h987f; 10'h131: x = 16'h97de; 10'h132: x = 16'h973c; 10'h133: x = 16'h9699; 10'h134: x = 16'h95f6; 10'h135: x = 16'h9553; 10'h136: x = 16'h94b0; 10'h137: x = 16'h940c; 10'h138: x = 16'h9368; 10'h139: x = 16'h92c3; 10'h13a: x = 16'h921e; 10'h13b: x = 16'h9179; 10'h13c: x = 16'h90d3; 10'h13d: x = 16'h902d; 10'h13e: x = 16'h8f87; 10'h13f: x = 16'h8ee0; 10'h140: x = 16'h8e39; 10'h141: x = 16'h8d92; 10'h142: x = 16'h8cea; 10'h143: x = 16'h8c42; 10'h144: x = 16'h8b9a; 10'h145: x = 16'h8af1; 10'h146: x = 16'h8a48; 10'h147: x = 16'h899f; 10'h148: x = 16'h88f5; 10'h149: x = 16'h884b; 10'h14a: x = 16'h87a1; 10'h14b: x = 16'h86f6; 10'h14c: x = 16'h864b; 10'h14d: x = 16'h85a0; 10'h14e: x = 16'h84f4; 10'h14f: x = 16'h8448; 10'h150: x = 16'h839c; 10'h151: x = 16'h82ef; 10'h152: x = 16'h8242; 10'h153: x = 16'h8195; 10'h154: x = 16'h80e7; 10'h155: x = 16'h803a; 10'h156: x = 16'h7f8b; 10'h157: x = 16'h7edd; 10'h158: x = 16'h7e2e; 10'h159: x = 16'h7d7f; 10'h15a: x = 16'h7cd0; 10'h15b: x = 16'h7c20; 10'h15c: x = 16'h7b70; 10'h15d: x = 16'h7ac0; 10'h15e: x = 16'h7a0f; 10'h15f: x = 16'h795e; 10'h160: x = 16'h78ad; 10'h161: x = 16'h77fb; 10'h162: x = 16'h774a; 10'h163: x = 16'h7698; 10'h164: x = 16'h75e5; 10'h165: x = 16'h7533; 10'h166: x = 16'h7480; 10'h167: x = 16'h73cd; 10'h168: x = 16'h7319; 10'h169: x = 16'h7265; 10'h16a: x = 16'h71b1; 10'h16b: x = 16'h70fd; 10'h16c: x = 16'h7049; 10'h16d: x = 16'h6f94; 10'h16e: x = 16'h6edf; 10'h16f: x = 16'h6e29; 10'h170: x = 16'h6d74; 10'h171: x = 16'h6cbe; 10'h172: x = 16'h6c08; 10'h173: x = 16'h6b51; 10'h174: x = 16'h6a9b; 10'h175: x = 16'h69e4; 10'h176: x = 16'h692d; 10'h177: x = 16'h6875; 10'h178: x = 16'h67bd; 10'h179: x = 16'h6705; 10'h17a: x = 16'h664d; 10'h17b: x = 16'h6595; 10'h17c: x = 16'h64dc; 10'h17d: x = 16'h6423; 10'h17e: x = 16'h636a; 10'h17f: x = 16'h62b1; 10'h180: x = 16'h61f7; 10'h181: x = 16'h613d; 10'h182: x = 16'h6083; 10'h183: x = 16'h5fc9; 10'h184: x = 16'h5f0e; 10'h185: x = 16'h5e53; 10'h186: x = 16'h5d98; 10'h187: x = 16'h5cdd; 10'h188: x = 16'h5c22; 10'h189: x = 16'h5b66; 10'h18a: x = 16'h5aaa; 10'h18b: x = 16'h59ee; 10'h18c: x = 16'h5931; 10'h18d: x = 16'h5875; 10'h18e: x = 16'h57b8; 10'h18f: x = 16'h56fb; 10'h190: x = 16'h563e; 10'h191: x = 16'h5581; 10'h192: x = 16'h54c3; 10'h193: x = 16'h5405; 10'h194: x = 16'h5347; 10'h195: x = 16'h5289; 10'h196: x = 16'h51ca; 10'h197: x = 16'h510c; 10'h198: x = 16'h504d; 10'h199: x = 16'h4f8e; 10'h19a: x = 16'h4ecf; 10'h19b: x = 16'h4e0f; 10'h19c: x = 16'h4d50; 10'h19d: x = 16'h4c90; 10'h19e: x = 16'h4bd0; 10'h19f: x = 16'h4b10; 10'h1a0: x = 16'h4a50; 10'h1a1: x = 16'h498f; 10'h1a2: x = 16'h48ce; 10'h1a3: x = 16'h480e; 10'h1a4: x = 16'h474d; 10'h1a5: x = 16'h468b; 10'h1a6: x = 16'h45ca; 10'h1a7: x = 16'h4508; 10'h1a8: x = 16'h4447; 10'h1a9: x = 16'h4385; 10'h1aa: x = 16'h42c3; 10'h1ab: x = 16'h4201; 10'h1ac: x = 16'h413e; 10'h1ad: x = 16'h407c; 10'h1ae: x = 16'h3fb9; 10'h1af: x = 16'h3ef6; 10'h1b0: x = 16'h3e33; 10'h1b1: x = 16'h3d70; 10'h1b2: x = 16'h3cad; 10'h1b3: x = 16'h3bea; 10'h1b4: x = 16'h3b26; 10'h1b5: x = 16'h3a62; 10'h1b6: x = 16'h399f; 10'h1b7: x = 16'h38db; 10'h1b8: x = 16'h3817; 10'h1b9: x = 16'h3752; 10'h1ba: x = 16'h368e; 10'h1bb: x = 16'h35c9; 10'h1bc: x = 16'h3505; 10'h1bd: x = 16'h3440; 10'h1be: x = 16'h337b; 10'h1bf: x = 16'h32b6; 10'h1c0: x = 16'h31f1; 10'h1c1: x = 16'h312c; 10'h1c2: x = 16'h3066; 10'h1c3: x = 16'h2fa1; 10'h1c4: x = 16'h2edb; 10'h1c5: x = 16'h2e15; 10'h1c6: x = 16'h2d50; 10'h1c7: x = 16'h2c8a; 10'h1c8: x = 16'h2bc4; 10'h1c9: x = 16'h2afe; 10'h1ca: x = 16'h2a37; 10'h1cb: x = 16'h2971; 10'h1cc: x = 16'h28aa; 10'h1cd: x = 16'h27e4; 10'h1ce: x = 16'h271d; 10'h1cf: x = 16'h2656; 10'h1d0: x = 16'h2590; 10'h1d1: x = 16'h24c9; 10'h1d2: x = 16'h2402; 10'h1d3: x = 16'h233b; 10'h1d4: x = 16'h2273; 10'h1d5: x = 16'h21ac; 10'h1d6: x = 16'h20e5; 10'h1d7: x = 16'h201d; 10'h1d8: x = 16'h1f56; 10'h1d9: x = 16'h1e8e; 10'h1da: x = 16'h1dc7; 10'h1db: x = 16'h1cff; 10'h1dc: x = 16'h1c37; 10'h1dd: x = 16'h1b6f; 10'h1de: x = 16'h1aa7; 10'h1df: x = 16'h19df; 10'h1e0: x = 16'h1917; 10'h1e1: x = 16'h184f; 10'h1e2: x = 16'h1787; 10'h1e3: x = 16'h16bf; 10'h1e4: x = 16'h15f6; 10'h1e5: x = 16'h152e; 10'h1e6: x = 16'h1466; 10'h1e7: x = 16'h139d; 10'h1e8: x = 16'h12d5; 10'h1e9: x = 16'h120c; 10'h1ea: x = 16'h1144; 10'h1eb: x = 16'h107b; 10'h1ec: x = 16'h fb2; 10'h1ed: x = 16'h eea; 10'h1ee: x = 16'h e21; 10'h1ef: x = 16'h d58; 10'h1f0: x = 16'h c8f; 10'h1f1: x = 16'h bc6; 10'h1f2: x = 16'h afe; 10'h1f3: x = 16'h a35; 10'h1f4: x = 16'h 96c; 10'h1f5: x = 16'h 8a3; 10'h1f6: x = 16'h 7da; 10'h1f7: x = 16'h 711; 10'h1f8: x = 16'h 648; 10'h1f9: x = 16'h 57f; 10'h1fa: x = 16'h 4b6; 10'h1fb: x = 16'h 3ed; 10'h1fc: x = 16'h 324; 10'h1fd: x = 16'h 25b; 10'h1fe: x = 16'h 192; 10'h1ff: x = 16'h  c9; 10'h200: x = 16'h   0; 10'h201: x = 16'hffffff37; 10'h202: x = 16'hfffffe6e; 10'h203: x = 16'hfffffda5; 10'h204: x = 16'hfffffcdc; 10'h205: x = 16'hfffffc13; 10'h206: x = 16'hfffffb4a; 10'h207: x = 16'hfffffa81; 10'h208: x = 16'hfffff9b8; 10'h209: x = 16'hfffff8ef; 10'h20a: x = 16'hfffff826; 10'h20b: x = 16'hfffff75d; 10'h20c: x = 16'hfffff694; 10'h20d: x = 16'hfffff5cb; 10'h20e: x = 16'hfffff502; 10'h20f: x = 16'hfffff43a; 10'h210: x = 16'hfffff371; 10'h211: x = 16'hfffff2a8; 10'h212: x = 16'hfffff1df; 10'h213: x = 16'hfffff116; 10'h214: x = 16'hfffff04e; 10'h215: x = 16'hffffef85; 10'h216: x = 16'hffffeebc; 10'h217: x = 16'hffffedf4; 10'h218: x = 16'hffffed2b; 10'h219: x = 16'hffffec63; 10'h21a: x = 16'hffffeb9a; 10'h21b: x = 16'hffffead2; 10'h21c: x = 16'hffffea0a; 10'h21d: x = 16'hffffe941; 10'h21e: x = 16'hffffe879; 10'h21f: x = 16'hffffe7b1; 10'h220: x = 16'hffffe6e9; 10'h221: x = 16'hffffe621; 10'h222: x = 16'hffffe559; 10'h223: x = 16'hffffe491; 10'h224: x = 16'hffffe3c9; 10'h225: x = 16'hffffe301; 10'h226: x = 16'hffffe239; 10'h227: x = 16'hffffe172; 10'h228: x = 16'hffffe0aa; 10'h229: x = 16'hffffdfe3; 10'h22a: x = 16'hffffdf1b; 10'h22b: x = 16'hffffde54; 10'h22c: x = 16'hffffdd8d; 10'h22d: x = 16'hffffdcc5; 10'h22e: x = 16'hffffdbfe; 10'h22f: x = 16'hffffdb37; 10'h230: x = 16'hffffda70; 10'h231: x = 16'hffffd9aa; 10'h232: x = 16'hffffd8e3; 10'h233: x = 16'hffffd81c; 10'h234: x = 16'hffffd756; 10'h235: x = 16'hffffd68f; 10'h236: x = 16'hffffd5c9; 10'h237: x = 16'hffffd502; 10'h238: x = 16'hffffd43c; 10'h239: x = 16'hffffd376; 10'h23a: x = 16'hffffd2b0; 10'h23b: x = 16'hffffd1eb; 10'h23c: x = 16'hffffd125; 10'h23d: x = 16'hffffd05f; 10'h23e: x = 16'hffffcf9a; 10'h23f: x = 16'hffffced4; 10'h240: x = 16'hffffce0f; 10'h241: x = 16'hffffcd4a; 10'h242: x = 16'hffffcc85; 10'h243: x = 16'hffffcbc0; 10'h244: x = 16'hffffcafb; 10'h245: x = 16'hffffca37; 10'h246: x = 16'hffffc972; 10'h247: x = 16'hffffc8ae; 10'h248: x = 16'hffffc7e9; 10'h249: x = 16'hffffc725; 10'h24a: x = 16'hffffc661; 10'h24b: x = 16'hffffc59e; 10'h24c: x = 16'hffffc4da; 10'h24d: x = 16'hffffc416; 10'h24e: x = 16'hffffc353; 10'h24f: x = 16'hffffc290; 10'h250: x = 16'hffffc1cd; 10'h251: x = 16'hffffc10a; 10'h252: x = 16'hffffc047; 10'h253: x = 16'hffffbf84; 10'h254: x = 16'hffffbec2; 10'h255: x = 16'hffffbdff; 10'h256: x = 16'hffffbd3d; 10'h257: x = 16'hffffbc7b; 10'h258: x = 16'hffffbbb9; 10'h259: x = 16'hffffbaf8; 10'h25a: x = 16'hffffba36; 10'h25b: x = 16'hffffb975; 10'h25c: x = 16'hffffb8b3; 10'h25d: x = 16'hffffb7f2; 10'h25e: x = 16'hffffb732; 10'h25f: x = 16'hffffb671; 10'h260: x = 16'hffffb5b0; 10'h261: x = 16'hffffb4f0; 10'h262: x = 16'hffffb430; 10'h263: x = 16'hffffb370; 10'h264: x = 16'hffffb2b0; 10'h265: x = 16'hffffb1f1; 10'h266: x = 16'hffffb131; 10'h267: x = 16'hffffb072; 10'h268: x = 16'hffffafb3; 10'h269: x = 16'hffffaef4; 10'h26a: x = 16'hffffae36; 10'h26b: x = 16'hffffad77; 10'h26c: x = 16'hffffacb9; 10'h26d: x = 16'hffffabfb; 10'h26e: x = 16'hffffab3d; 10'h26f: x = 16'hffffaa7f; 10'h270: x = 16'hffffa9c2; 10'h271: x = 16'hffffa905; 10'h272: x = 16'hffffa848; 10'h273: x = 16'hffffa78b; 10'h274: x = 16'hffffa6cf; 10'h275: x = 16'hffffa612; 10'h276: x = 16'hffffa556; 10'h277: x = 16'hffffa49a; 10'h278: x = 16'hffffa3de; 10'h279: x = 16'hffffa323; 10'h27a: x = 16'hffffa268; 10'h27b: x = 16'hffffa1ad; 10'h27c: x = 16'hffffa0f2; 10'h27d: x = 16'hffffa037; 10'h27e: x = 16'hffff9f7d; 10'h27f: x = 16'hffff9ec3; 10'h280: x = 16'hffff9e09; 10'h281: x = 16'hffff9d4f; 10'h282: x = 16'hffff9c96; 10'h283: x = 16'hffff9bdd; 10'h284: x = 16'hffff9b24; 10'h285: x = 16'hffff9a6b; 10'h286: x = 16'hffff99b3; 10'h287: x = 16'hffff98fb; 10'h288: x = 16'hffff9843; 10'h289: x = 16'hffff978b; 10'h28a: x = 16'hffff96d3; 10'h28b: x = 16'hffff961c; 10'h28c: x = 16'hffff9565; 10'h28d: x = 16'hffff94af; 10'h28e: x = 16'hffff93f8; 10'h28f: x = 16'hffff9342; 10'h290: x = 16'hffff928c; 10'h291: x = 16'hffff91d7; 10'h292: x = 16'hffff9121; 10'h293: x = 16'hffff906c; 10'h294: x = 16'hffff8fb7; 10'h295: x = 16'hffff8f03; 10'h296: x = 16'hffff8e4f; 10'h297: x = 16'hffff8d9b; 10'h298: x = 16'hffff8ce7; 10'h299: x = 16'hffff8c33; 10'h29a: x = 16'hffff8b80; 10'h29b: x = 16'hffff8acd; 10'h29c: x = 16'hffff8a1b; 10'h29d: x = 16'hffff8968; 10'h29e: x = 16'hffff88b6; 10'h29f: x = 16'hffff8805; 10'h2a0: x = 16'hffff8753; 10'h2a1: x = 16'hffff86a2; 10'h2a2: x = 16'hffff85f1; 10'h2a3: x = 16'hffff8540; 10'h2a4: x = 16'hffff8490; 10'h2a5: x = 16'hffff83e0; 10'h2a6: x = 16'hffff8330; 10'h2a7: x = 16'hffff8281; 10'h2a8: x = 16'hffff81d2; 10'h2a9: x = 16'hffff8123; 10'h2aa: x = 16'hffff8075; 10'h2ab: x = 16'hffff7fc6; 10'h2ac: x = 16'hffff7f19; 10'h2ad: x = 16'hffff7e6b; 10'h2ae: x = 16'hffff7dbe; 10'h2af: x = 16'hffff7d11; 10'h2b0: x = 16'hffff7c64; 10'h2b1: x = 16'hffff7bb8; 10'h2b2: x = 16'hffff7b0c; 10'h2b3: x = 16'hffff7a60; 10'h2b4: x = 16'hffff79b5; 10'h2b5: x = 16'hffff790a; 10'h2b6: x = 16'hffff785f; 10'h2b7: x = 16'hffff77b5; 10'h2b8: x = 16'hffff770b; 10'h2b9: x = 16'hffff7661; 10'h2ba: x = 16'hffff75b8; 10'h2bb: x = 16'hffff750f; 10'h2bc: x = 16'hffff7466; 10'h2bd: x = 16'hffff73be; 10'h2be: x = 16'hffff7316; 10'h2bf: x = 16'hffff726e; 10'h2c0: x = 16'hffff71c7; 10'h2c1: x = 16'hffff7120; 10'h2c2: x = 16'hffff7079; 10'h2c3: x = 16'hffff6fd3; 10'h2c4: x = 16'hffff6f2d; 10'h2c5: x = 16'hffff6e87; 10'h2c6: x = 16'hffff6de2; 10'h2c7: x = 16'hffff6d3d; 10'h2c8: x = 16'hffff6c98; 10'h2c9: x = 16'hffff6bf4; 10'h2ca: x = 16'hffff6b50; 10'h2cb: x = 16'hffff6aad; 10'h2cc: x = 16'hffff6a0a; 10'h2cd: x = 16'hffff6967; 10'h2ce: x = 16'hffff68c4; 10'h2cf: x = 16'hffff6822; 10'h2d0: x = 16'hffff6781; 10'h2d1: x = 16'hffff66df; 10'h2d2: x = 16'hffff663e; 10'h2d3: x = 16'hffff659e; 10'h2d4: x = 16'hffff64fe; 10'h2d5: x = 16'hffff645e; 10'h2d6: x = 16'hffff63be; 10'h2d7: x = 16'hffff631f; 10'h2d8: x = 16'hffff6281; 10'h2d9: x = 16'hffff61e2; 10'h2da: x = 16'hffff6144; 10'h2db: x = 16'hffff60a7; 10'h2dc: x = 16'hffff600a; 10'h2dd: x = 16'hffff5f6d; 10'h2de: x = 16'hffff5ed1; 10'h2df: x = 16'hffff5e35; 10'h2e0: x = 16'hffff5d99; 10'h2e1: x = 16'hffff5cfe; 10'h2e2: x = 16'hffff5c63; 10'h2e3: x = 16'hffff5bc8; 10'h2e4: x = 16'hffff5b2e; 10'h2e5: x = 16'hffff5a95; 10'h2e6: x = 16'hffff59fb; 10'h2e7: x = 16'hffff5963; 10'h2e8: x = 16'hffff58ca; 10'h2e9: x = 16'hffff5832; 10'h2ea: x = 16'hffff579a; 10'h2eb: x = 16'hffff5703; 10'h2ec: x = 16'hffff566c; 10'h2ed: x = 16'hffff55d6; 10'h2ee: x = 16'hffff5540; 10'h2ef: x = 16'hffff54aa; 10'h2f0: x = 16'hffff5415; 10'h2f1: x = 16'hffff5380; 10'h2f2: x = 16'hffff52ec; 10'h2f3: x = 16'hffff5258; 10'h2f4: x = 16'hffff51c5; 10'h2f5: x = 16'hffff5132; 10'h2f6: x = 16'hffff509f; 10'h2f7: x = 16'hffff500d; 10'h2f8: x = 16'hffff4f7b; 10'h2f9: x = 16'hffff4ee9; 10'h2fa: x = 16'hffff4e58; 10'h2fb: x = 16'hffff4dc8; 10'h2fc: x = 16'hffff4d38; 10'h2fd: x = 16'hffff4ca8; 10'h2fe: x = 16'hffff4c19; 10'h2ff: x = 16'hffff4b8a; 10'h300: x = 16'hffff4afc; 10'h301: x = 16'hffff4a6e; 10'h302: x = 16'hffff49e0; 10'h303: x = 16'hffff4953; 10'h304: x = 16'hffff48c6; 10'h305: x = 16'hffff483a; 10'h306: x = 16'hffff47ae; 10'h307: x = 16'hffff4723; 10'h308: x = 16'hffff4698; 10'h309: x = 16'hffff460e; 10'h30a: x = 16'hffff4584; 10'h30b: x = 16'hffff44fa; 10'h30c: x = 16'hffff4471; 10'h30d: x = 16'hffff43e9; 10'h30e: x = 16'hffff4360; 10'h30f: x = 16'hffff42d9; 10'h310: x = 16'hffff4252; 10'h311: x = 16'hffff41cb; 10'h312: x = 16'hffff4144; 10'h313: x = 16'hffff40bf; 10'h314: x = 16'hffff4039; 10'h315: x = 16'hffff3fb4; 10'h316: x = 16'hffff3f30; 10'h317: x = 16'hffff3eac; 10'h318: x = 16'hffff3e28; 10'h319: x = 16'hffff3da5; 10'h31a: x = 16'hffff3d22; 10'h31b: x = 16'hffff3ca0; 10'h31c: x = 16'hffff3c1e; 10'h31d: x = 16'hffff3b9d; 10'h31e: x = 16'hffff3b1d; 10'h31f: x = 16'hffff3a9c; 10'h320: x = 16'hffff3a1c; 10'h321: x = 16'hffff399d; 10'h322: x = 16'hffff391e; 10'h323: x = 16'hffff38a0; 10'h324: x = 16'hffff3822; 10'h325: x = 16'hffff37a5; 10'h326: x = 16'hffff3728; 10'h327: x = 16'hffff36ab; 10'h328: x = 16'hffff362f; 10'h329: x = 16'hffff35b4; 10'h32a: x = 16'hffff3539; 10'h32b: x = 16'hffff34bf; 10'h32c: x = 16'hffff3445; 10'h32d: x = 16'hffff33cb; 10'h32e: x = 16'hffff3352; 10'h32f: x = 16'hffff32da; 10'h330: x = 16'hffff3261; 10'h331: x = 16'hffff31ea; 10'h332: x = 16'hffff3173; 10'h333: x = 16'hffff30fc; 10'h334: x = 16'hffff3086; 10'h335: x = 16'hffff3011; 10'h336: x = 16'hffff2f9c; 10'h337: x = 16'hffff2f27; 10'h338: x = 16'hffff2eb3; 10'h339: x = 16'hffff2e40; 10'h33a: x = 16'hffff2dcd; 10'h33b: x = 16'hffff2d5a; 10'h33c: x = 16'hffff2ce8; 10'h33d: x = 16'hffff2c77; 10'h33e: x = 16'hffff2c06; 10'h33f: x = 16'hffff2b95; 10'h340: x = 16'hffff2b25; 10'h341: x = 16'hffff2ab6; 10'h342: x = 16'hffff2a47; 10'h343: x = 16'hffff29d9; 10'h344: x = 16'hffff296b; 10'h345: x = 16'hffff28fd; 10'h346: x = 16'hffff2890; 10'h347: x = 16'hffff2824; 10'h348: x = 16'hffff27b8; 10'h349: x = 16'hffff274d; 10'h34a: x = 16'hffff26e2; 10'h34b: x = 16'hffff2678; 10'h34c: x = 16'hffff260e; 10'h34d: x = 16'hffff25a5; 10'h34e: x = 16'hffff253c; 10'h34f: x = 16'hffff24d4; 10'h350: x = 16'hffff246c; 10'h351: x = 16'hffff2405; 10'h352: x = 16'hffff239f; 10'h353: x = 16'hffff2339; 10'h354: x = 16'hffff22d3; 10'h355: x = 16'hffff226e; 10'h356: x = 16'hffff220a; 10'h357: x = 16'hffff21a6; 10'h358: x = 16'hffff2142; 10'h359: x = 16'hffff20e0; 10'h35a: x = 16'hffff207d; 10'h35b: x = 16'hffff201c; 10'h35c: x = 16'hffff1fba; 10'h35d: x = 16'hffff1f5a; 10'h35e: x = 16'hffff1efa; 10'h35f: x = 16'hffff1e9a; 10'h360: x = 16'hffff1e3b; 10'h361: x = 16'hffff1ddc; 10'h362: x = 16'hffff1d7e; 10'h363: x = 16'hffff1d21; 10'h364: x = 16'hffff1cc4; 10'h365: x = 16'hffff1c68; 10'h366: x = 16'hffff1c0c; 10'h367: x = 16'hffff1bb1; 10'h368: x = 16'hffff1b56; 10'h369: x = 16'hffff1afc; 10'h36a: x = 16'hffff1aa2; 10'h36b: x = 16'hffff1a49; 10'h36c: x = 16'hffff19f1; 10'h36d: x = 16'hffff1999; 10'h36e: x = 16'hffff1942; 10'h36f: x = 16'hffff18eb; 10'h370: x = 16'hffff1895; 10'h371: x = 16'hffff183f; 10'h372: x = 16'hffff17ea; 10'h373: x = 16'hffff1795; 10'h374: x = 16'hffff1741; 10'h375: x = 16'hffff16ee; 10'h376: x = 16'hffff169b; 10'h377: x = 16'hffff1649; 10'h378: x = 16'hffff15f7; 10'h379: x = 16'hffff15a6; 10'h37a: x = 16'hffff1555; 10'h37b: x = 16'hffff1505; 10'h37c: x = 16'hffff14b5; 10'h37d: x = 16'hffff1467; 10'h37e: x = 16'hffff1418; 10'h37f: x = 16'hffff13ca; 10'h380: x = 16'hffff137d; 10'h381: x = 16'hffff1330; 10'h382: x = 16'hffff12e4; 10'h383: x = 16'hffff1299; 10'h384: x = 16'hffff124e; 10'h385: x = 16'hffff1204; 10'h386: x = 16'hffff11ba; 10'h387: x = 16'hffff1171; 10'h388: x = 16'hffff1128; 10'h389: x = 16'hffff10e0; 10'h38a: x = 16'hffff1098; 10'h38b: x = 16'hffff1051; 10'h38c: x = 16'hffff100b; 10'h38d: x = 16'hffff0fc5; 10'h38e: x = 16'hffff0f80; 10'h38f: x = 16'hffff0f3b; 10'h390: x = 16'hffff0ef7; 10'h391: x = 16'hffff0eb4; 10'h392: x = 16'hffff0e71; 10'h393: x = 16'hffff0e2f; 10'h394: x = 16'hffff0ded; 10'h395: x = 16'hffff0dac; 10'h396: x = 16'hffff0d6c; 10'h397: x = 16'hffff0d2c; 10'h398: x = 16'hffff0cec; 10'h399: x = 16'hffff0cad; 10'h39a: x = 16'hffff0c6f; 10'h39b: x = 16'hffff0c32; 10'h39c: x = 16'hffff0bf5; 10'h39d: x = 16'hffff0bb8; 10'h39e: x = 16'hffff0b7c; 10'h39f: x = 16'hffff0b41; 10'h3a0: x = 16'hffff0b06; 10'h3a1: x = 16'hffff0acc; 10'h3a2: x = 16'hffff0a93; 10'h3a3: x = 16'hffff0a5a; 10'h3a4: x = 16'hffff0a22; 10'h3a5: x = 16'hffff09ea; 10'h3a6: x = 16'hffff09b3; 10'h3a7: x = 16'hffff097c; 10'h3a8: x = 16'hffff0946; 10'h3a9: x = 16'hffff0911; 10'h3aa: x = 16'hffff08dc; 10'h3ab: x = 16'hffff08a8; 10'h3ac: x = 16'hffff0875; 10'h3ad: x = 16'hffff0842; 10'h3ae: x = 16'hffff080f; 10'h3af: x = 16'hffff07de; 10'h3b0: x = 16'hffff07ad; 10'h3b1: x = 16'hffff077c; 10'h3b2: x = 16'hffff074c; 10'h3b3: x = 16'hffff071d; 10'h3b4: x = 16'hffff06ee; 10'h3b5: x = 16'hffff06c0; 10'h3b6: x = 16'hffff0692; 10'h3b7: x = 16'hffff0665; 10'h3b8: x = 16'hffff0639; 10'h3b9: x = 16'hffff060d; 10'h3ba: x = 16'hffff05e2; 10'h3bb: x = 16'hffff05b7; 10'h3bc: x = 16'hffff058d; 10'h3bd: x = 16'hffff0564; 10'h3be: x = 16'hffff053b; 10'h3bf: x = 16'hffff0513; 10'h3c0: x = 16'hffff04ec; 10'h3c1: x = 16'hffff04c5; 10'h3c2: x = 16'hffff049f; 10'h3c3: x = 16'hffff0479; 10'h3c4: x = 16'hffff0454; 10'h3c5: x = 16'hffff042f; 10'h3c6: x = 16'hffff040b; 10'h3c7: x = 16'hffff03e8; 10'h3c8: x = 16'hffff03c5; 10'h3c9: x = 16'hffff03a3; 10'h3ca: x = 16'hffff0382; 10'h3cb: x = 16'hffff0361; 10'h3cc: x = 16'hffff0341; 10'h3cd: x = 16'hffff0321; 10'h3ce: x = 16'hffff0302; 10'h3cf: x = 16'hffff02e4; 10'h3d0: x = 16'hffff02c6; 10'h3d1: x = 16'hffff02a9; 10'h3d2: x = 16'hffff028c; 10'h3d3: x = 16'hffff0270; 10'h3d4: x = 16'hffff0255; 10'h3d5: x = 16'hffff023a; 10'h3d6: x = 16'hffff0220; 10'h3d7: x = 16'hffff0206; 10'h3d8: x = 16'hffff01ed; 10'h3d9: x = 16'hffff01d5; 10'h3da: x = 16'hffff01bd; 10'h3db: x = 16'hffff01a6; 10'h3dc: x = 16'hffff0190; 10'h3dd: x = 16'hffff017a; 10'h3de: x = 16'hffff0165; 10'h3df: x = 16'hffff0150; 10'h3e0: x = 16'hffff013c; 10'h3e1: x = 16'hffff0129; 10'h3e2: x = 16'hffff0116; 10'h3e3: x = 16'hffff0104; 10'h3e4: x = 16'hffff00f2; 10'h3e5: x = 16'hffff00e1; 10'h3e6: x = 16'hffff00d1; 10'h3e7: x = 16'hffff00c1; 10'h3e8: x = 16'hffff00b2; 10'h3e9: x = 16'hffff00a4; 10'h3ea: x = 16'hffff0096; 10'h3eb: x = 16'hffff0088; 10'h3ec: x = 16'hffff007c; 10'h3ed: x = 16'hffff0070; 10'h3ee: x = 16'hffff0064; 10'h3ef: x = 16'hffff005a; 10'h3f0: x = 16'hffff004f; 10'h3f1: x = 16'hffff0046; 10'h3f2: x = 16'hffff003d; 10'h3f3: x = 16'hffff0035; 10'h3f4: x = 16'hffff002d; 10'h3f5: x = 16'hffff0026; 10'h3f6: x = 16'hffff001f; 10'h3f7: x = 16'hffff0019; 10'h3f8: x = 16'hffff0014; 10'h3f9: x = 16'hffff0010; 10'h3fa: x = 16'hffff000c; 10'h3fb: x = 16'hffff0008; 10'h3fc: x = 16'hffff0005; 10'h3fd: x = 16'hffff0003; 10'h3fe: x = 16'hffff0002; 10'h3ff: x = 16'hffff0001; 			
		endcase
	end
endmodule

module sqrt_log (
	input	[11:0] data_in,
	output [15:0] data_out
);
	reg [15:0] x = 32'b0000_0000_0000_0000_0000_0000_0000_0000;
	
	assign data_out = x;
	
	always @(*) begin
		case(data_in)
		12'h  1: x = 16'h8284; 12'h  2: x = 16'h7cf5; 12'h  3: x = 16'h7997; 12'h  4: x = 16'h7725; 12'h  5: x = 16'h7536; 12'h  6: x = 16'h739b; 12'h  7: x = 16'h723c; 12'h  8: x = 16'h7108; 12'h  9: x = 16'h6ff5; 12'h  a: x = 16'h6efd; 12'h  b: x = 16'h6e1b; 12'h  c: x = 16'h6d4b; 12'h  d: x = 16'h6c8b; 12'h  e: x = 16'h6bd7; 12'h  f: x = 16'h6b2f; 12'h 10: x = 16'h6a91; 12'h 11: x = 16'h69fb; 12'h 12: x = 16'h696d; 12'h 13: x = 16'h68e7; 12'h 14: x = 16'h6866; 12'h 15: x = 16'h67eb; 12'h 16: x = 16'h6776; 12'h 17: x = 16'h6705; 12'h 18: x = 16'h6698; 12'h 19: x = 16'h6630; 12'h 1a: x = 16'h65cb; 12'h 1b: x = 16'h656a; 12'h 1c: x = 16'h650b; 12'h 1d: x = 16'h64b0; 12'h 1e: x = 16'h6458; 12'h 1f: x = 16'h6402; 12'h 20: x = 16'h63af; 12'h 21: x = 16'h635e; 12'h 22: x = 16'h630f; 12'h 23: x = 16'h62c2; 12'h 24: x = 16'h6277; 12'h 25: x = 16'h622e; 12'h 26: x = 16'h61e7; 12'h 27: x = 16'h61a1; 12'h 28: x = 16'h615d; 12'h 29: x = 16'h611a; 12'h 2a: x = 16'h60d9; 12'h 2b: x = 16'h6099; 12'h 2c: x = 16'h605b; 12'h 2d: x = 16'h601e; 12'h 2e: x = 16'h5fe2; 12'h 2f: x = 16'h5fa7; 12'h 30: x = 16'h5f6d; 12'h 31: x = 16'h5f34; 12'h 32: x = 16'h5efd; 12'h 33: x = 16'h5ec6; 12'h 34: x = 16'h5e90; 12'h 35: x = 16'h5e5b; 12'h 36: x = 16'h5e27; 12'h 37: x = 16'h5df4; 12'h 38: x = 16'h5dc2; 12'h 39: x = 16'h5d90; 12'h 3a: x = 16'h5d60; 12'h 3b: x = 16'h5d30; 12'h 3c: x = 16'h5d00; 12'h 3d: x = 16'h5cd2; 12'h 3e: x = 16'h5ca4; 12'h 3f: x = 16'h5c76; 12'h 40: x = 16'h5c4a; 12'h 41: x = 16'h5c1e; 12'h 42: x = 16'h5bf2; 12'h 43: x = 16'h5bc7; 12'h 44: x = 16'h5b9d; 12'h 45: x = 16'h5b73; 12'h 46: x = 16'h5b4a; 12'h 47: x = 16'h5b21; 12'h 48: x = 16'h5af9; 12'h 49: x = 16'h5ad1; 12'h 4a: x = 16'h5aaa; 12'h 4b: x = 16'h5a83; 12'h 4c: x = 16'h5a5c; 12'h 4d: x = 16'h5a36; 12'h 4e: x = 16'h5a11; 12'h 4f: x = 16'h59ec; 12'h 50: x = 16'h59c7; 12'h 51: x = 16'h59a3; 12'h 52: x = 16'h597f; 12'h 53: x = 16'h595b; 12'h 54: x = 16'h5938; 12'h 55: x = 16'h5915; 12'h 56: x = 16'h58f3; 12'h 57: x = 16'h58d1; 12'h 58: x = 16'h58af; 12'h 59: x = 16'h588e; 12'h 5a: x = 16'h586d; 12'h 5b: x = 16'h584c; 12'h 5c: x = 16'h582b; 12'h 5d: x = 16'h580b; 12'h 5e: x = 16'h57eb; 12'h 5f: x = 16'h57cc; 12'h 60: x = 16'h57ac; 12'h 61: x = 16'h578d; 12'h 62: x = 16'h576f; 12'h 63: x = 16'h5750; 12'h 64: x = 16'h5732; 12'h 65: x = 16'h5714; 12'h 66: x = 16'h56f6; 12'h 67: x = 16'h56d9; 12'h 68: x = 16'h56bc; 12'h 69: x = 16'h569f; 12'h 6a: x = 16'h5682; 12'h 6b: x = 16'h5666; 12'h 6c: x = 16'h5649; 12'h 6d: x = 16'h562d; 12'h 6e: x = 16'h5612; 12'h 6f: x = 16'h55f6; 12'h 70: x = 16'h55db; 12'h 71: x = 16'h55c0; 12'h 72: x = 16'h55a5; 12'h 73: x = 16'h558a; 12'h 74: x = 16'h556f; 12'h 75: x = 16'h5555; 12'h 76: x = 16'h553b; 12'h 77: x = 16'h5521; 12'h 78: x = 16'h5507; 12'h 79: x = 16'h54ed; 12'h 7a: x = 16'h54d4; 12'h 7b: x = 16'h54bb; 12'h 7c: x = 16'h54a2; 12'h 7d: x = 16'h5489; 12'h 7e: x = 16'h5470; 12'h 7f: x = 16'h5458; 12'h 80: x = 16'h543f; 12'h 81: x = 16'h5427; 12'h 82: x = 16'h540f; 12'h 83: x = 16'h53f7; 12'h 84: x = 16'h53df; 12'h 85: x = 16'h53c8; 12'h 86: x = 16'h53b0; 12'h 87: x = 16'h5399; 12'h 88: x = 16'h5382; 12'h 89: x = 16'h536b; 12'h 8a: x = 16'h5354; 12'h 8b: x = 16'h533d; 12'h 8c: x = 16'h5326; 12'h 8d: x = 16'h5310; 12'h 8e: x = 16'h52fa; 12'h 8f: x = 16'h52e4; 12'h 90: x = 16'h52cd; 12'h 91: x = 16'h52b8; 12'h 92: x = 16'h52a2; 12'h 93: x = 16'h528c; 12'h 94: x = 16'h5277; 12'h 95: x = 16'h5261; 12'h 96: x = 16'h524c; 12'h 97: x = 16'h5237; 12'h 98: x = 16'h5222; 12'h 99: x = 16'h520d; 12'h 9a: x = 16'h51f8; 12'h 9b: x = 16'h51e3; 12'h 9c: x = 16'h51cf; 12'h 9d: x = 16'h51ba; 12'h 9e: x = 16'h51a6; 12'h 9f: x = 16'h5191; 12'h a0: x = 16'h517d; 12'h a1: x = 16'h5169; 12'h a2: x = 16'h5155; 12'h a3: x = 16'h5141; 12'h a4: x = 16'h512e; 12'h a5: x = 16'h511a; 12'h a6: x = 16'h5107; 12'h a7: x = 16'h50f3; 12'h a8: x = 16'h50e0; 12'h a9: x = 16'h50cc; 12'h aa: x = 16'h50b9; 12'h ab: x = 16'h50a6; 12'h ac: x = 16'h5093; 12'h ad: x = 16'h5080; 12'h ae: x = 16'h506e; 12'h af: x = 16'h505b; 12'h b0: x = 16'h5048; 12'h b1: x = 16'h5036; 12'h b2: x = 16'h5023; 12'h b3: x = 16'h5011; 12'h b4: x = 16'h4fff; 12'h b5: x = 16'h4fed; 12'h b6: x = 16'h4fdb; 12'h b7: x = 16'h4fc9; 12'h b8: x = 16'h4fb7; 12'h b9: x = 16'h4fa5; 12'h ba: x = 16'h4f93; 12'h bb: x = 16'h4f81; 12'h bc: x = 16'h4f70; 12'h bd: x = 16'h4f5e; 12'h be: x = 16'h4f4d; 12'h bf: x = 16'h4f3c; 12'h c0: x = 16'h4f2a; 12'h c1: x = 16'h4f19; 12'h c2: x = 16'h4f08; 12'h c3: x = 16'h4ef7; 12'h c4: x = 16'h4ee6; 12'h c5: x = 16'h4ed5; 12'h c6: x = 16'h4ec4; 12'h c7: x = 16'h4eb3; 12'h c8: x = 16'h4ea3; 12'h c9: x = 16'h4e92; 12'h ca: x = 16'h4e81; 12'h cb: x = 16'h4e71; 12'h cc: x = 16'h4e61; 12'h cd: x = 16'h4e50; 12'h ce: x = 16'h4e40; 12'h cf: x = 16'h4e30; 12'h d0: x = 16'h4e1f; 12'h d1: x = 16'h4e0f; 12'h d2: x = 16'h4dff; 12'h d3: x = 16'h4def; 12'h d4: x = 16'h4ddf; 12'h d5: x = 16'h4dd0; 12'h d6: x = 16'h4dc0; 12'h d7: x = 16'h4db0; 12'h d8: x = 16'h4da0; 12'h d9: x = 16'h4d91; 12'h da: x = 16'h4d81; 12'h db: x = 16'h4d72; 12'h dc: x = 16'h4d62; 12'h dd: x = 16'h4d53; 12'h de: x = 16'h4d44; 12'h df: x = 16'h4d34; 12'h e0: x = 16'h4d25; 12'h e1: x = 16'h4d16; 12'h e2: x = 16'h4d07; 12'h e3: x = 16'h4cf8; 12'h e4: x = 16'h4ce9; 12'h e5: x = 16'h4cda; 12'h e6: x = 16'h4ccb; 12'h e7: x = 16'h4cbc; 12'h e8: x = 16'h4cae; 12'h e9: x = 16'h4c9f; 12'h ea: x = 16'h4c90; 12'h eb: x = 16'h4c82; 12'h ec: x = 16'h4c73; 12'h ed: x = 16'h4c65; 12'h ee: x = 16'h4c56; 12'h ef: x = 16'h4c48; 12'h f0: x = 16'h4c39; 12'h f1: x = 16'h4c2b; 12'h f2: x = 16'h4c1d; 12'h f3: x = 16'h4c0f; 12'h f4: x = 16'h4c00; 12'h f5: x = 16'h4bf2; 12'h f6: x = 16'h4be4; 12'h f7: x = 16'h4bd6; 12'h f8: x = 16'h4bc8; 12'h f9: x = 16'h4bba; 12'h fa: x = 16'h4bad; 12'h fb: x = 16'h4b9f; 12'h fc: x = 16'h4b91; 12'h fd: x = 16'h4b83; 12'h fe: x = 16'h4b75; 12'h ff: x = 16'h4b68; 12'h100: x = 16'h4b5a; 12'h101: x = 16'h4b4d; 12'h102: x = 16'h4b3f; 12'h103: x = 16'h4b32; 12'h104: x = 16'h4b24; 12'h105: x = 16'h4b17; 12'h106: x = 16'h4b09; 12'h107: x = 16'h4afc; 12'h108: x = 16'h4aef; 12'h109: x = 16'h4ae2; 12'h10a: x = 16'h4ad4; 12'h10b: x = 16'h4ac7; 12'h10c: x = 16'h4aba; 12'h10d: x = 16'h4aad; 12'h10e: x = 16'h4aa0; 12'h10f: x = 16'h4a93; 12'h110: x = 16'h4a86; 12'h111: x = 16'h4a79; 12'h112: x = 16'h4a6c; 12'h113: x = 16'h4a5f; 12'h114: x = 16'h4a53; 12'h115: x = 16'h4a46; 12'h116: x = 16'h4a39; 12'h117: x = 16'h4a2d; 12'h118: x = 16'h4a20; 12'h119: x = 16'h4a13; 12'h11a: x = 16'h4a07; 12'h11b: x = 16'h49fa; 12'h11c: x = 16'h49ee; 12'h11d: x = 16'h49e1; 12'h11e: x = 16'h49d5; 12'h11f: x = 16'h49c8; 12'h120: x = 16'h49bc; 12'h121: x = 16'h49b0; 12'h122: x = 16'h49a3; 12'h123: x = 16'h4997; 12'h124: x = 16'h498b; 12'h125: x = 16'h497f; 12'h126: x = 16'h4973; 12'h127: x = 16'h4966; 12'h128: x = 16'h495a; 12'h129: x = 16'h494e; 12'h12a: x = 16'h4942; 12'h12b: x = 16'h4936; 12'h12c: x = 16'h492a; 12'h12d: x = 16'h491e; 12'h12e: x = 16'h4912; 12'h12f: x = 16'h4907; 12'h130: x = 16'h48fb; 12'h131: x = 16'h48ef; 12'h132: x = 16'h48e3; 12'h133: x = 16'h48d7; 12'h134: x = 16'h48cc; 12'h135: x = 16'h48c0; 12'h136: x = 16'h48b4; 12'h137: x = 16'h48a9; 12'h138: x = 16'h489d; 12'h139: x = 16'h4892; 12'h13a: x = 16'h4886; 12'h13b: x = 16'h487b; 12'h13c: x = 16'h486f; 12'h13d: x = 16'h4864; 12'h13e: x = 16'h4858; 12'h13f: x = 16'h484d; 12'h140: x = 16'h4842; 12'h141: x = 16'h4836; 12'h142: x = 16'h482b; 12'h143: x = 16'h4820; 12'h144: x = 16'h4815; 12'h145: x = 16'h4809; 12'h146: x = 16'h47fe; 12'h147: x = 16'h47f3; 12'h148: x = 16'h47e8; 12'h149: x = 16'h47dd; 12'h14a: x = 16'h47d2; 12'h14b: x = 16'h47c7; 12'h14c: x = 16'h47bc; 12'h14d: x = 16'h47b1; 12'h14e: x = 16'h47a6; 12'h14f: x = 16'h479b; 12'h150: x = 16'h4790; 12'h151: x = 16'h4785; 12'h152: x = 16'h477a; 12'h153: x = 16'h476f; 12'h154: x = 16'h4764; 12'h155: x = 16'h475a; 12'h156: x = 16'h474f; 12'h157: x = 16'h4744; 12'h158: x = 16'h4739; 12'h159: x = 16'h472f; 12'h15a: x = 16'h4724; 12'h15b: x = 16'h4719; 12'h15c: x = 16'h470f; 12'h15d: x = 16'h4704; 12'h15e: x = 16'h46fa; 12'h15f: x = 16'h46ef; 12'h160: x = 16'h46e5; 12'h161: x = 16'h46da; 12'h162: x = 16'h46d0; 12'h163: x = 16'h46c5; 12'h164: x = 16'h46bb; 12'h165: x = 16'h46b0; 12'h166: x = 16'h46a6; 12'h167: x = 16'h469c; 12'h168: x = 16'h4691; 12'h169: x = 16'h4687; 12'h16a: x = 16'h467d; 12'h16b: x = 16'h4672; 12'h16c: x = 16'h4668; 12'h16d: x = 16'h465e; 12'h16e: x = 16'h4654; 12'h16f: x = 16'h464a; 12'h170: x = 16'h463f; 12'h171: x = 16'h4635; 12'h172: x = 16'h462b; 12'h173: x = 16'h4621; 12'h174: x = 16'h4617; 12'h175: x = 16'h460d; 12'h176: x = 16'h4603; 12'h177: x = 16'h45f9; 12'h178: x = 16'h45ef; 12'h179: x = 16'h45e5; 12'h17a: x = 16'h45db; 12'h17b: x = 16'h45d1; 12'h17c: x = 16'h45c7; 12'h17d: x = 16'h45bd; 12'h17e: x = 16'h45b4; 12'h17f: x = 16'h45aa; 12'h180: x = 16'h45a0; 12'h181: x = 16'h4596; 12'h182: x = 16'h458c; 12'h183: x = 16'h4583; 12'h184: x = 16'h4579; 12'h185: x = 16'h456f; 12'h186: x = 16'h4565; 12'h187: x = 16'h455c; 12'h188: x = 16'h4552; 12'h189: x = 16'h4548; 12'h18a: x = 16'h453f; 12'h18b: x = 16'h4535; 12'h18c: x = 16'h452c; 12'h18d: x = 16'h4522; 12'h18e: x = 16'h4519; 12'h18f: x = 16'h450f; 12'h190: x = 16'h4506; 12'h191: x = 16'h44fc; 12'h192: x = 16'h44f3; 12'h193: x = 16'h44e9; 12'h194: x = 16'h44e0; 12'h195: x = 16'h44d6; 12'h196: x = 16'h44cd; 12'h197: x = 16'h44c4; 12'h198: x = 16'h44ba; 12'h199: x = 16'h44b1; 12'h19a: x = 16'h44a8; 12'h19b: x = 16'h449e; 12'h19c: x = 16'h4495; 12'h19d: x = 16'h448c; 12'h19e: x = 16'h4482; 12'h19f: x = 16'h4479; 12'h1a0: x = 16'h4470; 12'h1a1: x = 16'h4467; 12'h1a2: x = 16'h445e; 12'h1a3: x = 16'h4454; 12'h1a4: x = 16'h444b; 12'h1a5: x = 16'h4442; 12'h1a6: x = 16'h4439; 12'h1a7: x = 16'h4430; 12'h1a8: x = 16'h4427; 12'h1a9: x = 16'h441e; 12'h1aa: x = 16'h4415; 12'h1ab: x = 16'h440c; 12'h1ac: x = 16'h4403; 12'h1ad: x = 16'h43fa; 12'h1ae: x = 16'h43f1; 12'h1af: x = 16'h43e8; 12'h1b0: x = 16'h43df; 12'h1b1: x = 16'h43d6; 12'h1b2: x = 16'h43cd; 12'h1b3: x = 16'h43c4; 12'h1b4: x = 16'h43bb; 12'h1b5: x = 16'h43b2; 12'h1b6: x = 16'h43a9; 12'h1b7: x = 16'h43a1; 12'h1b8: x = 16'h4398; 12'h1b9: x = 16'h438f; 12'h1ba: x = 16'h4386; 12'h1bb: x = 16'h437d; 12'h1bc: x = 16'h4375; 12'h1bd: x = 16'h436c; 12'h1be: x = 16'h4363; 12'h1bf: x = 16'h435a; 12'h1c0: x = 16'h4352; 12'h1c1: x = 16'h4349; 12'h1c2: x = 16'h4340; 12'h1c3: x = 16'h4338; 12'h1c4: x = 16'h432f; 12'h1c5: x = 16'h4327; 12'h1c6: x = 16'h431e; 12'h1c7: x = 16'h4315; 12'h1c8: x = 16'h430d; 12'h1c9: x = 16'h4304; 12'h1ca: x = 16'h42fc; 12'h1cb: x = 16'h42f3; 12'h1cc: x = 16'h42eb; 12'h1cd: x = 16'h42e2; 12'h1ce: x = 16'h42da; 12'h1cf: x = 16'h42d1; 12'h1d0: x = 16'h42c9; 12'h1d1: x = 16'h42c0; 12'h1d2: x = 16'h42b8; 12'h1d3: x = 16'h42af; 12'h1d4: x = 16'h42a7; 12'h1d5: x = 16'h429e; 12'h1d6: x = 16'h4296; 12'h1d7: x = 16'h428e; 12'h1d8: x = 16'h4285; 12'h1d9: x = 16'h427d; 12'h1da: x = 16'h4275; 12'h1db: x = 16'h426c; 12'h1dc: x = 16'h4264; 12'h1dd: x = 16'h425c; 12'h1de: x = 16'h4254; 12'h1df: x = 16'h424b; 12'h1e0: x = 16'h4243; 12'h1e1: x = 16'h423b; 12'h1e2: x = 16'h4233; 12'h1e3: x = 16'h422a; 12'h1e4: x = 16'h4222; 12'h1e5: x = 16'h421a; 12'h1e6: x = 16'h4212; 12'h1e7: x = 16'h420a; 12'h1e8: x = 16'h4201; 12'h1e9: x = 16'h41f9; 12'h1ea: x = 16'h41f1; 12'h1eb: x = 16'h41e9; 12'h1ec: x = 16'h41e1; 12'h1ed: x = 16'h41d9; 12'h1ee: x = 16'h41d1; 12'h1ef: x = 16'h41c9; 12'h1f0: x = 16'h41c1; 12'h1f1: x = 16'h41b9; 12'h1f2: x = 16'h41b1; 12'h1f3: x = 16'h41a9; 12'h1f4: x = 16'h41a1; 12'h1f5: x = 16'h4199; 12'h1f6: x = 16'h4191; 12'h1f7: x = 16'h4189; 12'h1f8: x = 16'h4181; 12'h1f9: x = 16'h4179; 12'h1fa: x = 16'h4171; 12'h1fb: x = 16'h4169; 12'h1fc: x = 16'h4161; 12'h1fd: x = 16'h4159; 12'h1fe: x = 16'h4151; 12'h1ff: x = 16'h414a; 12'h200: x = 16'h4142; 12'h201: x = 16'h413a; 12'h202: x = 16'h4132; 12'h203: x = 16'h412a; 12'h204: x = 16'h4122; 12'h205: x = 16'h411b; 12'h206: x = 16'h4113; 12'h207: x = 16'h410b; 12'h208: x = 16'h4103; 12'h209: x = 16'h40fc; 12'h20a: x = 16'h40f4; 12'h20b: x = 16'h40ec; 12'h20c: x = 16'h40e4; 12'h20d: x = 16'h40dd; 12'h20e: x = 16'h40d5; 12'h20f: x = 16'h40cd; 12'h210: x = 16'h40c6; 12'h211: x = 16'h40be; 12'h212: x = 16'h40b6; 12'h213: x = 16'h40af; 12'h214: x = 16'h40a7; 12'h215: x = 16'h409f; 12'h216: x = 16'h4098; 12'h217: x = 16'h4090; 12'h218: x = 16'h4089; 12'h219: x = 16'h4081; 12'h21a: x = 16'h407a; 12'h21b: x = 16'h4072; 12'h21c: x = 16'h406a; 12'h21d: x = 16'h4063; 12'h21e: x = 16'h405b; 12'h21f: x = 16'h4054; 12'h220: x = 16'h404c; 12'h221: x = 16'h4045; 12'h222: x = 16'h403d; 12'h223: x = 16'h4036; 12'h224: x = 16'h402e; 12'h225: x = 16'h4027; 12'h226: x = 16'h4020; 12'h227: x = 16'h4018; 12'h228: x = 16'h4011; 12'h229: x = 16'h4009; 12'h22a: x = 16'h4002; 12'h22b: x = 16'h3ffb; 12'h22c: x = 16'h3ff3; 12'h22d: x = 16'h3fec; 12'h22e: x = 16'h3fe4; 12'h22f: x = 16'h3fdd; 12'h230: x = 16'h3fd6; 12'h231: x = 16'h3fce; 12'h232: x = 16'h3fc7; 12'h233: x = 16'h3fc0; 12'h234: x = 16'h3fb9; 12'h235: x = 16'h3fb1; 12'h236: x = 16'h3faa; 12'h237: x = 16'h3fa3; 12'h238: x = 16'h3f9b; 12'h239: x = 16'h3f94; 12'h23a: x = 16'h3f8d; 12'h23b: x = 16'h3f86; 12'h23c: x = 16'h3f7e; 12'h23d: x = 16'h3f77; 12'h23e: x = 16'h3f70; 12'h23f: x = 16'h3f69; 12'h240: x = 16'h3f62; 12'h241: x = 16'h3f5b; 12'h242: x = 16'h3f53; 12'h243: x = 16'h3f4c; 12'h244: x = 16'h3f45; 12'h245: x = 16'h3f3e; 12'h246: x = 16'h3f37; 12'h247: x = 16'h3f30; 12'h248: x = 16'h3f29; 12'h249: x = 16'h3f21; 12'h24a: x = 16'h3f1a; 12'h24b: x = 16'h3f13; 12'h24c: x = 16'h3f0c; 12'h24d: x = 16'h3f05; 12'h24e: x = 16'h3efe; 12'h24f: x = 16'h3ef7; 12'h250: x = 16'h3ef0; 12'h251: x = 16'h3ee9; 12'h252: x = 16'h3ee2; 12'h253: x = 16'h3edb; 12'h254: x = 16'h3ed4; 12'h255: x = 16'h3ecd; 12'h256: x = 16'h3ec6; 12'h257: x = 16'h3ebf; 12'h258: x = 16'h3eb8; 12'h259: x = 16'h3eb1; 12'h25a: x = 16'h3eaa; 12'h25b: x = 16'h3ea3; 12'h25c: x = 16'h3e9c; 12'h25d: x = 16'h3e95; 12'h25e: x = 16'h3e8e; 12'h25f: x = 16'h3e87; 12'h260: x = 16'h3e81; 12'h261: x = 16'h3e7a; 12'h262: x = 16'h3e73; 12'h263: x = 16'h3e6c; 12'h264: x = 16'h3e65; 12'h265: x = 16'h3e5e; 12'h266: x = 16'h3e57; 12'h267: x = 16'h3e50; 12'h268: x = 16'h3e4a; 12'h269: x = 16'h3e43; 12'h26a: x = 16'h3e3c; 12'h26b: x = 16'h3e35; 12'h26c: x = 16'h3e2e; 12'h26d: x = 16'h3e28; 12'h26e: x = 16'h3e21; 12'h26f: x = 16'h3e1a; 12'h270: x = 16'h3e13; 12'h271: x = 16'h3e0c; 12'h272: x = 16'h3e06; 12'h273: x = 16'h3dff; 12'h274: x = 16'h3df8; 12'h275: x = 16'h3df1; 12'h276: x = 16'h3deb; 12'h277: x = 16'h3de4; 12'h278: x = 16'h3ddd; 12'h279: x = 16'h3dd7; 12'h27a: x = 16'h3dd0; 12'h27b: x = 16'h3dc9; 12'h27c: x = 16'h3dc3; 12'h27d: x = 16'h3dbc; 12'h27e: x = 16'h3db5; 12'h27f: x = 16'h3daf; 12'h280: x = 16'h3da8; 12'h281: x = 16'h3da1; 12'h282: x = 16'h3d9b; 12'h283: x = 16'h3d94; 12'h284: x = 16'h3d8d; 12'h285: x = 16'h3d87; 12'h286: x = 16'h3d80; 12'h287: x = 16'h3d7a; 12'h288: x = 16'h3d73; 12'h289: x = 16'h3d6c; 12'h28a: x = 16'h3d66; 12'h28b: x = 16'h3d5f; 12'h28c: x = 16'h3d59; 12'h28d: x = 16'h3d52; 12'h28e: x = 16'h3d4c; 12'h28f: x = 16'h3d45; 12'h290: x = 16'h3d3f; 12'h291: x = 16'h3d38; 12'h292: x = 16'h3d32; 12'h293: x = 16'h3d2b; 12'h294: x = 16'h3d25; 12'h295: x = 16'h3d1e; 12'h296: x = 16'h3d18; 12'h297: x = 16'h3d11; 12'h298: x = 16'h3d0b; 12'h299: x = 16'h3d04; 12'h29a: x = 16'h3cfe; 12'h29b: x = 16'h3cf7; 12'h29c: x = 16'h3cf1; 12'h29d: x = 16'h3cea; 12'h29e: x = 16'h3ce4; 12'h29f: x = 16'h3cde; 12'h2a0: x = 16'h3cd7; 12'h2a1: x = 16'h3cd1; 12'h2a2: x = 16'h3cca; 12'h2a3: x = 16'h3cc4; 12'h2a4: x = 16'h3cbe; 12'h2a5: x = 16'h3cb7; 12'h2a6: x = 16'h3cb1; 12'h2a7: x = 16'h3caa; 12'h2a8: x = 16'h3ca4; 12'h2a9: x = 16'h3c9e; 12'h2aa: x = 16'h3c97; 12'h2ab: x = 16'h3c91; 12'h2ac: x = 16'h3c8b; 12'h2ad: x = 16'h3c84; 12'h2ae: x = 16'h3c7e; 12'h2af: x = 16'h3c78; 12'h2b0: x = 16'h3c71; 12'h2b1: x = 16'h3c6b; 12'h2b2: x = 16'h3c65; 12'h2b3: x = 16'h3c5f; 12'h2b4: x = 16'h3c58; 12'h2b5: x = 16'h3c52; 12'h2b6: x = 16'h3c4c; 12'h2b7: x = 16'h3c45; 12'h2b8: x = 16'h3c3f; 12'h2b9: x = 16'h3c39; 12'h2ba: x = 16'h3c33; 12'h2bb: x = 16'h3c2c; 12'h2bc: x = 16'h3c26; 12'h2bd: x = 16'h3c20; 12'h2be: x = 16'h3c1a; 12'h2bf: x = 16'h3c14; 12'h2c0: x = 16'h3c0d; 12'h2c1: x = 16'h3c07; 12'h2c2: x = 16'h3c01; 12'h2c3: x = 16'h3bfb; 12'h2c4: x = 16'h3bf5; 12'h2c5: x = 16'h3bee; 12'h2c6: x = 16'h3be8; 12'h2c7: x = 16'h3be2; 12'h2c8: x = 16'h3bdc; 12'h2c9: x = 16'h3bd6; 12'h2ca: x = 16'h3bd0; 12'h2cb: x = 16'h3bca; 12'h2cc: x = 16'h3bc3; 12'h2cd: x = 16'h3bbd; 12'h2ce: x = 16'h3bb7; 12'h2cf: x = 16'h3bb1; 12'h2d0: x = 16'h3bab; 12'h2d1: x = 16'h3ba5; 12'h2d2: x = 16'h3b9f; 12'h2d3: x = 16'h3b99; 12'h2d4: x = 16'h3b93; 12'h2d5: x = 16'h3b8d; 12'h2d6: x = 16'h3b86; 12'h2d7: x = 16'h3b80; 12'h2d8: x = 16'h3b7a; 12'h2d9: x = 16'h3b74; 12'h2da: x = 16'h3b6e; 12'h2db: x = 16'h3b68; 12'h2dc: x = 16'h3b62; 12'h2dd: x = 16'h3b5c; 12'h2de: x = 16'h3b56; 12'h2df: x = 16'h3b50; 12'h2e0: x = 16'h3b4a; 12'h2e1: x = 16'h3b44; 12'h2e2: x = 16'h3b3e; 12'h2e3: x = 16'h3b38; 12'h2e4: x = 16'h3b32; 12'h2e5: x = 16'h3b2c; 12'h2e6: x = 16'h3b26; 12'h2e7: x = 16'h3b20; 12'h2e8: x = 16'h3b1a; 12'h2e9: x = 16'h3b14; 12'h2ea: x = 16'h3b0e; 12'h2eb: x = 16'h3b08; 12'h2ec: x = 16'h3b02; 12'h2ed: x = 16'h3afc; 12'h2ee: x = 16'h3af7; 12'h2ef: x = 16'h3af1; 12'h2f0: x = 16'h3aeb; 12'h2f1: x = 16'h3ae5; 12'h2f2: x = 16'h3adf; 12'h2f3: x = 16'h3ad9; 12'h2f4: x = 16'h3ad3; 12'h2f5: x = 16'h3acd; 12'h2f6: x = 16'h3ac7; 12'h2f7: x = 16'h3ac1; 12'h2f8: x = 16'h3abc; 12'h2f9: x = 16'h3ab6; 12'h2fa: x = 16'h3ab0; 12'h2fb: x = 16'h3aaa; 12'h2fc: x = 16'h3aa4; 12'h2fd: x = 16'h3a9e; 12'h2fe: x = 16'h3a98; 12'h2ff: x = 16'h3a93; 12'h300: x = 16'h3a8d; 12'h301: x = 16'h3a87; 12'h302: x = 16'h3a81; 12'h303: x = 16'h3a7b; 12'h304: x = 16'h3a75; 12'h305: x = 16'h3a70; 12'h306: x = 16'h3a6a; 12'h307: x = 16'h3a64; 12'h308: x = 16'h3a5e; 12'h309: x = 16'h3a58; 12'h30a: x = 16'h3a53; 12'h30b: x = 16'h3a4d; 12'h30c: x = 16'h3a47; 12'h30d: x = 16'h3a41; 12'h30e: x = 16'h3a3c; 12'h30f: x = 16'h3a36; 12'h310: x = 16'h3a30; 12'h311: x = 16'h3a2a; 12'h312: x = 16'h3a25; 12'h313: x = 16'h3a1f; 12'h314: x = 16'h3a19; 12'h315: x = 16'h3a13; 12'h316: x = 16'h3a0e; 12'h317: x = 16'h3a08; 12'h318: x = 16'h3a02; 12'h319: x = 16'h39fd; 12'h31a: x = 16'h39f7; 12'h31b: x = 16'h39f1; 12'h31c: x = 16'h39ec; 12'h31d: x = 16'h39e6; 12'h31e: x = 16'h39e0; 12'h31f: x = 16'h39db; 12'h320: x = 16'h39d5; 12'h321: x = 16'h39cf; 12'h322: x = 16'h39ca; 12'h323: x = 16'h39c4; 12'h324: x = 16'h39be; 12'h325: x = 16'h39b9; 12'h326: x = 16'h39b3; 12'h327: x = 16'h39ad; 12'h328: x = 16'h39a8; 12'h329: x = 16'h39a2; 12'h32a: x = 16'h399c; 12'h32b: x = 16'h3997; 12'h32c: x = 16'h3991; 12'h32d: x = 16'h398c; 12'h32e: x = 16'h3986; 12'h32f: x = 16'h3980; 12'h330: x = 16'h397b; 12'h331: x = 16'h3975; 12'h332: x = 16'h3970; 12'h333: x = 16'h396a; 12'h334: x = 16'h3964; 12'h335: x = 16'h395f; 12'h336: x = 16'h3959; 12'h337: x = 16'h3954; 12'h338: x = 16'h394e; 12'h339: x = 16'h3949; 12'h33a: x = 16'h3943; 12'h33b: x = 16'h393e; 12'h33c: x = 16'h3938; 12'h33d: x = 16'h3933; 12'h33e: x = 16'h392d; 12'h33f: x = 16'h3928; 12'h340: x = 16'h3922; 12'h341: x = 16'h391c; 12'h342: x = 16'h3917; 12'h343: x = 16'h3911; 12'h344: x = 16'h390c; 12'h345: x = 16'h3906; 12'h346: x = 16'h3901; 12'h347: x = 16'h38fb; 12'h348: x = 16'h38f6; 12'h349: x = 16'h38f1; 12'h34a: x = 16'h38eb; 12'h34b: x = 16'h38e6; 12'h34c: x = 16'h38e0; 12'h34d: x = 16'h38db; 12'h34e: x = 16'h38d5; 12'h34f: x = 16'h38d0; 12'h350: x = 16'h38ca; 12'h351: x = 16'h38c5; 12'h352: x = 16'h38bf; 12'h353: x = 16'h38ba; 12'h354: x = 16'h38b5; 12'h355: x = 16'h38af; 12'h356: x = 16'h38aa; 12'h357: x = 16'h38a4; 12'h358: x = 16'h389f; 12'h359: x = 16'h389a; 12'h35a: x = 16'h3894; 12'h35b: x = 16'h388f; 12'h35c: x = 16'h3889; 12'h35d: x = 16'h3884; 12'h35e: x = 16'h387f; 12'h35f: x = 16'h3879; 12'h360: x = 16'h3874; 12'h361: x = 16'h386e; 12'h362: x = 16'h3869; 12'h363: x = 16'h3864; 12'h364: x = 16'h385e; 12'h365: x = 16'h3859; 12'h366: x = 16'h3854; 12'h367: x = 16'h384e; 12'h368: x = 16'h3849; 12'h369: x = 16'h3844; 12'h36a: x = 16'h383e; 12'h36b: x = 16'h3839; 12'h36c: x = 16'h3834; 12'h36d: x = 16'h382e; 12'h36e: x = 16'h3829; 12'h36f: x = 16'h3824; 12'h370: x = 16'h381e; 12'h371: x = 16'h3819; 12'h372: x = 16'h3814; 12'h373: x = 16'h380e; 12'h374: x = 16'h3809; 12'h375: x = 16'h3804; 12'h376: x = 16'h37ff; 12'h377: x = 16'h37f9; 12'h378: x = 16'h37f4; 12'h379: x = 16'h37ef; 12'h37a: x = 16'h37e9; 12'h37b: x = 16'h37e4; 12'h37c: x = 16'h37df; 12'h37d: x = 16'h37da; 12'h37e: x = 16'h37d4; 12'h37f: x = 16'h37cf; 12'h380: x = 16'h37ca; 12'h381: x = 16'h37c5; 12'h382: x = 16'h37bf; 12'h383: x = 16'h37ba; 12'h384: x = 16'h37b5; 12'h385: x = 16'h37b0; 12'h386: x = 16'h37ab; 12'h387: x = 16'h37a5; 12'h388: x = 16'h37a0; 12'h389: x = 16'h379b; 12'h38a: x = 16'h3796; 12'h38b: x = 16'h3790; 12'h38c: x = 16'h378b; 12'h38d: x = 16'h3786; 12'h38e: x = 16'h3781; 12'h38f: x = 16'h377c; 12'h390: x = 16'h3777; 12'h391: x = 16'h3771; 12'h392: x = 16'h376c; 12'h393: x = 16'h3767; 12'h394: x = 16'h3762; 12'h395: x = 16'h375d; 12'h396: x = 16'h3757; 12'h397: x = 16'h3752; 12'h398: x = 16'h374d; 12'h399: x = 16'h3748; 12'h39a: x = 16'h3743; 12'h39b: x = 16'h373e; 12'h39c: x = 16'h3739; 12'h39d: x = 16'h3733; 12'h39e: x = 16'h372e; 12'h39f: x = 16'h3729; 12'h3a0: x = 16'h3724; 12'h3a1: x = 16'h371f; 12'h3a2: x = 16'h371a; 12'h3a3: x = 16'h3715; 12'h3a4: x = 16'h3710; 12'h3a5: x = 16'h370b; 12'h3a6: x = 16'h3705; 12'h3a7: x = 16'h3700; 12'h3a8: x = 16'h36fb; 12'h3a9: x = 16'h36f6; 12'h3aa: x = 16'h36f1; 12'h3ab: x = 16'h36ec; 12'h3ac: x = 16'h36e7; 12'h3ad: x = 16'h36e2; 12'h3ae: x = 16'h36dd; 12'h3af: x = 16'h36d8; 12'h3b0: x = 16'h36d3; 12'h3b1: x = 16'h36ce; 12'h3b2: x = 16'h36c8; 12'h3b3: x = 16'h36c3; 12'h3b4: x = 16'h36be; 12'h3b5: x = 16'h36b9; 12'h3b6: x = 16'h36b4; 12'h3b7: x = 16'h36af; 12'h3b8: x = 16'h36aa; 12'h3b9: x = 16'h36a5; 12'h3ba: x = 16'h36a0; 12'h3bb: x = 16'h369b; 12'h3bc: x = 16'h3696; 12'h3bd: x = 16'h3691; 12'h3be: x = 16'h368c; 12'h3bf: x = 16'h3687; 12'h3c0: x = 16'h3682; 12'h3c1: x = 16'h367d; 12'h3c2: x = 16'h3678; 12'h3c3: x = 16'h3673; 12'h3c4: x = 16'h366e; 12'h3c5: x = 16'h3669; 12'h3c6: x = 16'h3664; 12'h3c7: x = 16'h365f; 12'h3c8: x = 16'h365a; 12'h3c9: x = 16'h3655; 12'h3ca: x = 16'h3650; 12'h3cb: x = 16'h364b; 12'h3cc: x = 16'h3646; 12'h3cd: x = 16'h3641; 12'h3ce: x = 16'h363c; 12'h3cf: x = 16'h3637; 12'h3d0: x = 16'h3632; 12'h3d1: x = 16'h362d; 12'h3d2: x = 16'h3628; 12'h3d3: x = 16'h3623; 12'h3d4: x = 16'h361e; 12'h3d5: x = 16'h361a; 12'h3d6: x = 16'h3615; 12'h3d7: x = 16'h3610; 12'h3d8: x = 16'h360b; 12'h3d9: x = 16'h3606; 12'h3da: x = 16'h3601; 12'h3db: x = 16'h35fc; 12'h3dc: x = 16'h35f7; 12'h3dd: x = 16'h35f2; 12'h3de: x = 16'h35ed; 12'h3df: x = 16'h35e8; 12'h3e0: x = 16'h35e3; 12'h3e1: x = 16'h35de; 12'h3e2: x = 16'h35da; 12'h3e3: x = 16'h35d5; 12'h3e4: x = 16'h35d0; 12'h3e5: x = 16'h35cb; 12'h3e6: x = 16'h35c6; 12'h3e7: x = 16'h35c1; 12'h3e8: x = 16'h35bc; 12'h3e9: x = 16'h35b7; 12'h3ea: x = 16'h35b3; 12'h3eb: x = 16'h35ae; 12'h3ec: x = 16'h35a9; 12'h3ed: x = 16'h35a4; 12'h3ee: x = 16'h359f; 12'h3ef: x = 16'h359a; 12'h3f0: x = 16'h3595; 12'h3f1: x = 16'h3590; 12'h3f2: x = 16'h358c; 12'h3f3: x = 16'h3587; 12'h3f4: x = 16'h3582; 12'h3f5: x = 16'h357d; 12'h3f6: x = 16'h3578; 12'h3f7: x = 16'h3573; 12'h3f8: x = 16'h356f; 12'h3f9: x = 16'h356a; 12'h3fa: x = 16'h3565; 12'h3fb: x = 16'h3560; 12'h3fc: x = 16'h355b; 12'h3fd: x = 16'h3557; 12'h3fe: x = 16'h3552; 12'h3ff: x = 16'h354d; 12'h400: x = 16'h3548; 12'h401: x = 16'h3543; 12'h402: x = 16'h353e; 12'h403: x = 16'h353a; 12'h404: x = 16'h3535; 12'h405: x = 16'h3530; 12'h406: x = 16'h352b; 12'h407: x = 16'h3527; 12'h408: x = 16'h3522; 12'h409: x = 16'h351d; 12'h40a: x = 16'h3518; 12'h40b: x = 16'h3513; 12'h40c: x = 16'h350f; 12'h40d: x = 16'h350a; 12'h40e: x = 16'h3505; 12'h40f: x = 16'h3500; 12'h410: x = 16'h34fc; 12'h411: x = 16'h34f7; 12'h412: x = 16'h34f2; 12'h413: x = 16'h34ed; 12'h414: x = 16'h34e9; 12'h415: x = 16'h34e4; 12'h416: x = 16'h34df; 12'h417: x = 16'h34da; 12'h418: x = 16'h34d6; 12'h419: x = 16'h34d1; 12'h41a: x = 16'h34cc; 12'h41b: x = 16'h34c7; 12'h41c: x = 16'h34c3; 12'h41d: x = 16'h34be; 12'h41e: x = 16'h34b9; 12'h41f: x = 16'h34b5; 12'h420: x = 16'h34b0; 12'h421: x = 16'h34ab; 12'h422: x = 16'h34a6; 12'h423: x = 16'h34a2; 12'h424: x = 16'h349d; 12'h425: x = 16'h3498; 12'h426: x = 16'h3494; 12'h427: x = 16'h348f; 12'h428: x = 16'h348a; 12'h429: x = 16'h3486; 12'h42a: x = 16'h3481; 12'h42b: x = 16'h347c; 12'h42c: x = 16'h3477; 12'h42d: x = 16'h3473; 12'h42e: x = 16'h346e; 12'h42f: x = 16'h3469; 12'h430: x = 16'h3465; 12'h431: x = 16'h3460; 12'h432: x = 16'h345b; 12'h433: x = 16'h3457; 12'h434: x = 16'h3452; 12'h435: x = 16'h344e; 12'h436: x = 16'h3449; 12'h437: x = 16'h3444; 12'h438: x = 16'h3440; 12'h439: x = 16'h343b; 12'h43a: x = 16'h3436; 12'h43b: x = 16'h3432; 12'h43c: x = 16'h342d; 12'h43d: x = 16'h3428; 12'h43e: x = 16'h3424; 12'h43f: x = 16'h341f; 12'h440: x = 16'h341a; 12'h441: x = 16'h3416; 12'h442: x = 16'h3411; 12'h443: x = 16'h340d; 12'h444: x = 16'h3408; 12'h445: x = 16'h3403; 12'h446: x = 16'h33ff; 12'h447: x = 16'h33fa; 12'h448: x = 16'h33f6; 12'h449: x = 16'h33f1; 12'h44a: x = 16'h33ec; 12'h44b: x = 16'h33e8; 12'h44c: x = 16'h33e3; 12'h44d: x = 16'h33df; 12'h44e: x = 16'h33da; 12'h44f: x = 16'h33d5; 12'h450: x = 16'h33d1; 12'h451: x = 16'h33cc; 12'h452: x = 16'h33c8; 12'h453: x = 16'h33c3; 12'h454: x = 16'h33bf; 12'h455: x = 16'h33ba; 12'h456: x = 16'h33b5; 12'h457: x = 16'h33b1; 12'h458: x = 16'h33ac; 12'h459: x = 16'h33a8; 12'h45a: x = 16'h33a3; 12'h45b: x = 16'h339f; 12'h45c: x = 16'h339a; 12'h45d: x = 16'h3395; 12'h45e: x = 16'h3391; 12'h45f: x = 16'h338c; 12'h460: x = 16'h3388; 12'h461: x = 16'h3383; 12'h462: x = 16'h337f; 12'h463: x = 16'h337a; 12'h464: x = 16'h3376; 12'h465: x = 16'h3371; 12'h466: x = 16'h336d; 12'h467: x = 16'h3368; 12'h468: x = 16'h3364; 12'h469: x = 16'h335f; 12'h46a: x = 16'h335b; 12'h46b: x = 16'h3356; 12'h46c: x = 16'h3352; 12'h46d: x = 16'h334d; 12'h46e: x = 16'h3348; 12'h46f: x = 16'h3344; 12'h470: x = 16'h333f; 12'h471: x = 16'h333b; 12'h472: x = 16'h3336; 12'h473: x = 16'h3332; 12'h474: x = 16'h332d; 12'h475: x = 16'h3329; 12'h476: x = 16'h3325; 12'h477: x = 16'h3320; 12'h478: x = 16'h331c; 12'h479: x = 16'h3317; 12'h47a: x = 16'h3313; 12'h47b: x = 16'h330e; 12'h47c: x = 16'h330a; 12'h47d: x = 16'h3305; 12'h47e: x = 16'h3301; 12'h47f: x = 16'h32fc; 12'h480: x = 16'h32f8; 12'h481: x = 16'h32f3; 12'h482: x = 16'h32ef; 12'h483: x = 16'h32ea; 12'h484: x = 16'h32e6; 12'h485: x = 16'h32e1; 12'h486: x = 16'h32dd; 12'h487: x = 16'h32d9; 12'h488: x = 16'h32d4; 12'h489: x = 16'h32d0; 12'h48a: x = 16'h32cb; 12'h48b: x = 16'h32c7; 12'h48c: x = 16'h32c2; 12'h48d: x = 16'h32be; 12'h48e: x = 16'h32b9; 12'h48f: x = 16'h32b5; 12'h490: x = 16'h32b1; 12'h491: x = 16'h32ac; 12'h492: x = 16'h32a8; 12'h493: x = 16'h32a3; 12'h494: x = 16'h329f; 12'h495: x = 16'h329b; 12'h496: x = 16'h3296; 12'h497: x = 16'h3292; 12'h498: x = 16'h328d; 12'h499: x = 16'h3289; 12'h49a: x = 16'h3284; 12'h49b: x = 16'h3280; 12'h49c: x = 16'h327c; 12'h49d: x = 16'h3277; 12'h49e: x = 16'h3273; 12'h49f: x = 16'h326e; 12'h4a0: x = 16'h326a; 12'h4a1: x = 16'h3266; 12'h4a2: x = 16'h3261; 12'h4a3: x = 16'h325d; 12'h4a4: x = 16'h3259; 12'h4a5: x = 16'h3254; 12'h4a6: x = 16'h3250; 12'h4a7: x = 16'h324b; 12'h4a8: x = 16'h3247; 12'h4a9: x = 16'h3243; 12'h4aa: x = 16'h323e; 12'h4ab: x = 16'h323a; 12'h4ac: x = 16'h3236; 12'h4ad: x = 16'h3231; 12'h4ae: x = 16'h322d; 12'h4af: x = 16'h3228; 12'h4b0: x = 16'h3224; 12'h4b1: x = 16'h3220; 12'h4b2: x = 16'h321b; 12'h4b3: x = 16'h3217; 12'h4b4: x = 16'h3213; 12'h4b5: x = 16'h320e; 12'h4b6: x = 16'h320a; 12'h4b7: x = 16'h3206; 12'h4b8: x = 16'h3201; 12'h4b9: x = 16'h31fd; 12'h4ba: x = 16'h31f9; 12'h4bb: x = 16'h31f4; 12'h4bc: x = 16'h31f0; 12'h4bd: x = 16'h31ec; 12'h4be: x = 16'h31e7; 12'h4bf: x = 16'h31e3; 12'h4c0: x = 16'h31df; 12'h4c1: x = 16'h31da; 12'h4c2: x = 16'h31d6; 12'h4c3: x = 16'h31d2; 12'h4c4: x = 16'h31cd; 12'h4c5: x = 16'h31c9; 12'h4c6: x = 16'h31c5; 12'h4c7: x = 16'h31c0; 12'h4c8: x = 16'h31bc; 12'h4c9: x = 16'h31b8; 12'h4ca: x = 16'h31b4; 12'h4cb: x = 16'h31af; 12'h4cc: x = 16'h31ab; 12'h4cd: x = 16'h31a7; 12'h4ce: x = 16'h31a2; 12'h4cf: x = 16'h319e; 12'h4d0: x = 16'h319a; 12'h4d1: x = 16'h3195; 12'h4d2: x = 16'h3191; 12'h4d3: x = 16'h318d; 12'h4d4: x = 16'h3189; 12'h4d5: x = 16'h3184; 12'h4d6: x = 16'h3180; 12'h4d7: x = 16'h317c; 12'h4d8: x = 16'h3177; 12'h4d9: x = 16'h3173; 12'h4da: x = 16'h316f; 12'h4db: x = 16'h316b; 12'h4dc: x = 16'h3166; 12'h4dd: x = 16'h3162; 12'h4de: x = 16'h315e; 12'h4df: x = 16'h315a; 12'h4e0: x = 16'h3155; 12'h4e1: x = 16'h3151; 12'h4e2: x = 16'h314d; 12'h4e3: x = 16'h3149; 12'h4e4: x = 16'h3144; 12'h4e5: x = 16'h3140; 12'h4e6: x = 16'h313c; 12'h4e7: x = 16'h3138; 12'h4e8: x = 16'h3133; 12'h4e9: x = 16'h312f; 12'h4ea: x = 16'h312b; 12'h4eb: x = 16'h3127; 12'h4ec: x = 16'h3122; 12'h4ed: x = 16'h311e; 12'h4ee: x = 16'h311a; 12'h4ef: x = 16'h3116; 12'h4f0: x = 16'h3111; 12'h4f1: x = 16'h310d; 12'h4f2: x = 16'h3109; 12'h4f3: x = 16'h3105; 12'h4f4: x = 16'h3101; 12'h4f5: x = 16'h30fc; 12'h4f6: x = 16'h30f8; 12'h4f7: x = 16'h30f4; 12'h4f8: x = 16'h30f0; 12'h4f9: x = 16'h30ec; 12'h4fa: x = 16'h30e7; 12'h4fb: x = 16'h30e3; 12'h4fc: x = 16'h30df; 12'h4fd: x = 16'h30db; 12'h4fe: x = 16'h30d7; 12'h4ff: x = 16'h30d2; 12'h500: x = 16'h30ce; 12'h501: x = 16'h30ca; 12'h502: x = 16'h30c6; 12'h503: x = 16'h30c2; 12'h504: x = 16'h30bd; 12'h505: x = 16'h30b9; 12'h506: x = 16'h30b5; 12'h507: x = 16'h30b1; 12'h508: x = 16'h30ad; 12'h509: x = 16'h30a8; 12'h50a: x = 16'h30a4; 12'h50b: x = 16'h30a0; 12'h50c: x = 16'h309c; 12'h50d: x = 16'h3098; 12'h50e: x = 16'h3094; 12'h50f: x = 16'h308f; 12'h510: x = 16'h308b; 12'h511: x = 16'h3087; 12'h512: x = 16'h3083; 12'h513: x = 16'h307f; 12'h514: x = 16'h307b; 12'h515: x = 16'h3076; 12'h516: x = 16'h3072; 12'h517: x = 16'h306e; 12'h518: x = 16'h306a; 12'h519: x = 16'h3066; 12'h51a: x = 16'h3062; 12'h51b: x = 16'h305d; 12'h51c: x = 16'h3059; 12'h51d: x = 16'h3055; 12'h51e: x = 16'h3051; 12'h51f: x = 16'h304d; 12'h520: x = 16'h3049; 12'h521: x = 16'h3045; 12'h522: x = 16'h3041; 12'h523: x = 16'h303c; 12'h524: x = 16'h3038; 12'h525: x = 16'h3034; 12'h526: x = 16'h3030; 12'h527: x = 16'h302c; 12'h528: x = 16'h3028; 12'h529: x = 16'h3024; 12'h52a: x = 16'h301f; 12'h52b: x = 16'h301b; 12'h52c: x = 16'h3017; 12'h52d: x = 16'h3013; 12'h52e: x = 16'h300f; 12'h52f: x = 16'h300b; 12'h530: x = 16'h3007; 12'h531: x = 16'h3003; 12'h532: x = 16'h2fff; 12'h533: x = 16'h2ffa; 12'h534: x = 16'h2ff6; 12'h535: x = 16'h2ff2; 12'h536: x = 16'h2fee; 12'h537: x = 16'h2fea; 12'h538: x = 16'h2fe6; 12'h539: x = 16'h2fe2; 12'h53a: x = 16'h2fde; 12'h53b: x = 16'h2fda; 12'h53c: x = 16'h2fd6; 12'h53d: x = 16'h2fd2; 12'h53e: x = 16'h2fcd; 12'h53f: x = 16'h2fc9; 12'h540: x = 16'h2fc5; 12'h541: x = 16'h2fc1; 12'h542: x = 16'h2fbd; 12'h543: x = 16'h2fb9; 12'h544: x = 16'h2fb5; 12'h545: x = 16'h2fb1; 12'h546: x = 16'h2fad; 12'h547: x = 16'h2fa9; 12'h548: x = 16'h2fa5; 12'h549: x = 16'h2fa1; 12'h54a: x = 16'h2f9d; 12'h54b: x = 16'h2f98; 12'h54c: x = 16'h2f94; 12'h54d: x = 16'h2f90; 12'h54e: x = 16'h2f8c; 12'h54f: x = 16'h2f88; 12'h550: x = 16'h2f84; 12'h551: x = 16'h2f80; 12'h552: x = 16'h2f7c; 12'h553: x = 16'h2f78; 12'h554: x = 16'h2f74; 12'h555: x = 16'h2f70; 12'h556: x = 16'h2f6c; 12'h557: x = 16'h2f68; 12'h558: x = 16'h2f64; 12'h559: x = 16'h2f60; 12'h55a: x = 16'h2f5c; 12'h55b: x = 16'h2f58; 12'h55c: x = 16'h2f54; 12'h55d: x = 16'h2f50; 12'h55e: x = 16'h2f4c; 12'h55f: x = 16'h2f47; 12'h560: x = 16'h2f43; 12'h561: x = 16'h2f3f; 12'h562: x = 16'h2f3b; 12'h563: x = 16'h2f37; 12'h564: x = 16'h2f33; 12'h565: x = 16'h2f2f; 12'h566: x = 16'h2f2b; 12'h567: x = 16'h2f27; 12'h568: x = 16'h2f23; 12'h569: x = 16'h2f1f; 12'h56a: x = 16'h2f1b; 12'h56b: x = 16'h2f17; 12'h56c: x = 16'h2f13; 12'h56d: x = 16'h2f0f; 12'h56e: x = 16'h2f0b; 12'h56f: x = 16'h2f07; 12'h570: x = 16'h2f03; 12'h571: x = 16'h2eff; 12'h572: x = 16'h2efb; 12'h573: x = 16'h2ef7; 12'h574: x = 16'h2ef3; 12'h575: x = 16'h2eef; 12'h576: x = 16'h2eeb; 12'h577: x = 16'h2ee7; 12'h578: x = 16'h2ee3; 12'h579: x = 16'h2edf; 12'h57a: x = 16'h2edb; 12'h57b: x = 16'h2ed7; 12'h57c: x = 16'h2ed3; 12'h57d: x = 16'h2ecf; 12'h57e: x = 16'h2ecb; 12'h57f: x = 16'h2ec7; 12'h580: x = 16'h2ec3; 12'h581: x = 16'h2ebf; 12'h582: x = 16'h2ebb; 12'h583: x = 16'h2eb7; 12'h584: x = 16'h2eb3; 12'h585: x = 16'h2eaf; 12'h586: x = 16'h2eab; 12'h587: x = 16'h2ea7; 12'h588: x = 16'h2ea3; 12'h589: x = 16'h2e9f; 12'h58a: x = 16'h2e9c; 12'h58b: x = 16'h2e98; 12'h58c: x = 16'h2e94; 12'h58d: x = 16'h2e90; 12'h58e: x = 16'h2e8c; 12'h58f: x = 16'h2e88; 12'h590: x = 16'h2e84; 12'h591: x = 16'h2e80; 12'h592: x = 16'h2e7c; 12'h593: x = 16'h2e78; 12'h594: x = 16'h2e74; 12'h595: x = 16'h2e70; 12'h596: x = 16'h2e6c; 12'h597: x = 16'h2e68; 12'h598: x = 16'h2e64; 12'h599: x = 16'h2e60; 12'h59a: x = 16'h2e5c; 12'h59b: x = 16'h2e58; 12'h59c: x = 16'h2e54; 12'h59d: x = 16'h2e50; 12'h59e: x = 16'h2e4c; 12'h59f: x = 16'h2e49; 12'h5a0: x = 16'h2e45; 12'h5a1: x = 16'h2e41; 12'h5a2: x = 16'h2e3d; 12'h5a3: x = 16'h2e39; 12'h5a4: x = 16'h2e35; 12'h5a5: x = 16'h2e31; 12'h5a6: x = 16'h2e2d; 12'h5a7: x = 16'h2e29; 12'h5a8: x = 16'h2e25; 12'h5a9: x = 16'h2e21; 12'h5aa: x = 16'h2e1d; 12'h5ab: x = 16'h2e19; 12'h5ac: x = 16'h2e16; 12'h5ad: x = 16'h2e12; 12'h5ae: x = 16'h2e0e; 12'h5af: x = 16'h2e0a; 12'h5b0: x = 16'h2e06; 12'h5b1: x = 16'h2e02; 12'h5b2: x = 16'h2dfe; 12'h5b3: x = 16'h2dfa; 12'h5b4: x = 16'h2df6; 12'h5b5: x = 16'h2df2; 12'h5b6: x = 16'h2dee; 12'h5b7: x = 16'h2deb; 12'h5b8: x = 16'h2de7; 12'h5b9: x = 16'h2de3; 12'h5ba: x = 16'h2ddf; 12'h5bb: x = 16'h2ddb; 12'h5bc: x = 16'h2dd7; 12'h5bd: x = 16'h2dd3; 12'h5be: x = 16'h2dcf; 12'h5bf: x = 16'h2dcb; 12'h5c0: x = 16'h2dc7; 12'h5c1: x = 16'h2dc4; 12'h5c2: x = 16'h2dc0; 12'h5c3: x = 16'h2dbc; 12'h5c4: x = 16'h2db8; 12'h5c5: x = 16'h2db4; 12'h5c6: x = 16'h2db0; 12'h5c7: x = 16'h2dac; 12'h5c8: x = 16'h2da8; 12'h5c9: x = 16'h2da4; 12'h5ca: x = 16'h2da1; 12'h5cb: x = 16'h2d9d; 12'h5cc: x = 16'h2d99; 12'h5cd: x = 16'h2d95; 12'h5ce: x = 16'h2d91; 12'h5cf: x = 16'h2d8d; 12'h5d0: x = 16'h2d89; 12'h5d1: x = 16'h2d86; 12'h5d2: x = 16'h2d82; 12'h5d3: x = 16'h2d7e; 12'h5d4: x = 16'h2d7a; 12'h5d5: x = 16'h2d76; 12'h5d6: x = 16'h2d72; 12'h5d7: x = 16'h2d6e; 12'h5d8: x = 16'h2d6a; 12'h5d9: x = 16'h2d67; 12'h5da: x = 16'h2d63; 12'h5db: x = 16'h2d5f; 12'h5dc: x = 16'h2d5b; 12'h5dd: x = 16'h2d57; 12'h5de: x = 16'h2d53; 12'h5df: x = 16'h2d4f; 12'h5e0: x = 16'h2d4c; 12'h5e1: x = 16'h2d48; 12'h5e2: x = 16'h2d44; 12'h5e3: x = 16'h2d40; 12'h5e4: x = 16'h2d3c; 12'h5e5: x = 16'h2d38; 12'h5e6: x = 16'h2d35; 12'h5e7: x = 16'h2d31; 12'h5e8: x = 16'h2d2d; 12'h5e9: x = 16'h2d29; 12'h5ea: x = 16'h2d25; 12'h5eb: x = 16'h2d21; 12'h5ec: x = 16'h2d1e; 12'h5ed: x = 16'h2d1a; 12'h5ee: x = 16'h2d16; 12'h5ef: x = 16'h2d12; 12'h5f0: x = 16'h2d0e; 12'h5f1: x = 16'h2d0a; 12'h5f2: x = 16'h2d07; 12'h5f3: x = 16'h2d03; 12'h5f4: x = 16'h2cff; 12'h5f5: x = 16'h2cfb; 12'h5f6: x = 16'h2cf7; 12'h5f7: x = 16'h2cf3; 12'h5f8: x = 16'h2cf0; 12'h5f9: x = 16'h2cec; 12'h5fa: x = 16'h2ce8; 12'h5fb: x = 16'h2ce4; 12'h5fc: x = 16'h2ce0; 12'h5fd: x = 16'h2cdd; 12'h5fe: x = 16'h2cd9; 12'h5ff: x = 16'h2cd5; 12'h600: x = 16'h2cd1; 12'h601: x = 16'h2ccd; 12'h602: x = 16'h2cca; 12'h603: x = 16'h2cc6; 12'h604: x = 16'h2cc2; 12'h605: x = 16'h2cbe; 12'h606: x = 16'h2cba; 12'h607: x = 16'h2cb7; 12'h608: x = 16'h2cb3; 12'h609: x = 16'h2caf; 12'h60a: x = 16'h2cab; 12'h60b: x = 16'h2ca7; 12'h60c: x = 16'h2ca4; 12'h60d: x = 16'h2ca0; 12'h60e: x = 16'h2c9c; 12'h60f: x = 16'h2c98; 12'h610: x = 16'h2c94; 12'h611: x = 16'h2c91; 12'h612: x = 16'h2c8d; 12'h613: x = 16'h2c89; 12'h614: x = 16'h2c85; 12'h615: x = 16'h2c81; 12'h616: x = 16'h2c7e; 12'h617: x = 16'h2c7a; 12'h618: x = 16'h2c76; 12'h619: x = 16'h2c72; 12'h61a: x = 16'h2c6f; 12'h61b: x = 16'h2c6b; 12'h61c: x = 16'h2c67; 12'h61d: x = 16'h2c63; 12'h61e: x = 16'h2c5f; 12'h61f: x = 16'h2c5c; 12'h620: x = 16'h2c58; 12'h621: x = 16'h2c54; 12'h622: x = 16'h2c50; 12'h623: x = 16'h2c4d; 12'h624: x = 16'h2c49; 12'h625: x = 16'h2c45; 12'h626: x = 16'h2c41; 12'h627: x = 16'h2c3e; 12'h628: x = 16'h2c3a; 12'h629: x = 16'h2c36; 12'h62a: x = 16'h2c32; 12'h62b: x = 16'h2c2f; 12'h62c: x = 16'h2c2b; 12'h62d: x = 16'h2c27; 12'h62e: x = 16'h2c23; 12'h62f: x = 16'h2c1f; 12'h630: x = 16'h2c1c; 12'h631: x = 16'h2c18; 12'h632: x = 16'h2c14; 12'h633: x = 16'h2c10; 12'h634: x = 16'h2c0d; 12'h635: x = 16'h2c09; 12'h636: x = 16'h2c05; 12'h637: x = 16'h2c01; 12'h638: x = 16'h2bfe; 12'h639: x = 16'h2bfa; 12'h63a: x = 16'h2bf6; 12'h63b: x = 16'h2bf3; 12'h63c: x = 16'h2bef; 12'h63d: x = 16'h2beb; 12'h63e: x = 16'h2be7; 12'h63f: x = 16'h2be4; 12'h640: x = 16'h2be0; 12'h641: x = 16'h2bdc; 12'h642: x = 16'h2bd8; 12'h643: x = 16'h2bd5; 12'h644: x = 16'h2bd1; 12'h645: x = 16'h2bcd; 12'h646: x = 16'h2bc9; 12'h647: x = 16'h2bc6; 12'h648: x = 16'h2bc2; 12'h649: x = 16'h2bbe; 12'h64a: x = 16'h2bbb; 12'h64b: x = 16'h2bb7; 12'h64c: x = 16'h2bb3; 12'h64d: x = 16'h2baf; 12'h64e: x = 16'h2bac; 12'h64f: x = 16'h2ba8; 12'h650: x = 16'h2ba4; 12'h651: x = 16'h2ba1; 12'h652: x = 16'h2b9d; 12'h653: x = 16'h2b99; 12'h654: x = 16'h2b95; 12'h655: x = 16'h2b92; 12'h656: x = 16'h2b8e; 12'h657: x = 16'h2b8a; 12'h658: x = 16'h2b87; 12'h659: x = 16'h2b83; 12'h65a: x = 16'h2b7f; 12'h65b: x = 16'h2b7b; 12'h65c: x = 16'h2b78; 12'h65d: x = 16'h2b74; 12'h65e: x = 16'h2b70; 12'h65f: x = 16'h2b6d; 12'h660: x = 16'h2b69; 12'h661: x = 16'h2b65; 12'h662: x = 16'h2b62; 12'h663: x = 16'h2b5e; 12'h664: x = 16'h2b5a; 12'h665: x = 16'h2b56; 12'h666: x = 16'h2b53; 12'h667: x = 16'h2b4f; 12'h668: x = 16'h2b4b; 12'h669: x = 16'h2b48; 12'h66a: x = 16'h2b44; 12'h66b: x = 16'h2b40; 12'h66c: x = 16'h2b3d; 12'h66d: x = 16'h2b39; 12'h66e: x = 16'h2b35; 12'h66f: x = 16'h2b32; 12'h670: x = 16'h2b2e; 12'h671: x = 16'h2b2a; 12'h672: x = 16'h2b26; 12'h673: x = 16'h2b23; 12'h674: x = 16'h2b1f; 12'h675: x = 16'h2b1b; 12'h676: x = 16'h2b18; 12'h677: x = 16'h2b14; 12'h678: x = 16'h2b10; 12'h679: x = 16'h2b0d; 12'h67a: x = 16'h2b09; 12'h67b: x = 16'h2b05; 12'h67c: x = 16'h2b02; 12'h67d: x = 16'h2afe; 12'h67e: x = 16'h2afa; 12'h67f: x = 16'h2af7; 12'h680: x = 16'h2af3; 12'h681: x = 16'h2aef; 12'h682: x = 16'h2aec; 12'h683: x = 16'h2ae8; 12'h684: x = 16'h2ae4; 12'h685: x = 16'h2ae1; 12'h686: x = 16'h2add; 12'h687: x = 16'h2ad9; 12'h688: x = 16'h2ad6; 12'h689: x = 16'h2ad2; 12'h68a: x = 16'h2ace; 12'h68b: x = 16'h2acb; 12'h68c: x = 16'h2ac7; 12'h68d: x = 16'h2ac3; 12'h68e: x = 16'h2ac0; 12'h68f: x = 16'h2abc; 12'h690: x = 16'h2ab8; 12'h691: x = 16'h2ab5; 12'h692: x = 16'h2ab1; 12'h693: x = 16'h2aae; 12'h694: x = 16'h2aaa; 12'h695: x = 16'h2aa6; 12'h696: x = 16'h2aa3; 12'h697: x = 16'h2a9f; 12'h698: x = 16'h2a9b; 12'h699: x = 16'h2a98; 12'h69a: x = 16'h2a94; 12'h69b: x = 16'h2a90; 12'h69c: x = 16'h2a8d; 12'h69d: x = 16'h2a89; 12'h69e: x = 16'h2a85; 12'h69f: x = 16'h2a82; 12'h6a0: x = 16'h2a7e; 12'h6a1: x = 16'h2a7b; 12'h6a2: x = 16'h2a77; 12'h6a3: x = 16'h2a73; 12'h6a4: x = 16'h2a70; 12'h6a5: x = 16'h2a6c; 12'h6a6: x = 16'h2a68; 12'h6a7: x = 16'h2a65; 12'h6a8: x = 16'h2a61; 12'h6a9: x = 16'h2a5d; 12'h6aa: x = 16'h2a5a; 12'h6ab: x = 16'h2a56; 12'h6ac: x = 16'h2a53; 12'h6ad: x = 16'h2a4f; 12'h6ae: x = 16'h2a4b; 12'h6af: x = 16'h2a48; 12'h6b0: x = 16'h2a44; 12'h6b1: x = 16'h2a40; 12'h6b2: x = 16'h2a3d; 12'h6b3: x = 16'h2a39; 12'h6b4: x = 16'h2a36; 12'h6b5: x = 16'h2a32; 12'h6b6: x = 16'h2a2e; 12'h6b7: x = 16'h2a2b; 12'h6b8: x = 16'h2a27; 12'h6b9: x = 16'h2a23; 12'h6ba: x = 16'h2a20; 12'h6bb: x = 16'h2a1c; 12'h6bc: x = 16'h2a19; 12'h6bd: x = 16'h2a15; 12'h6be: x = 16'h2a11; 12'h6bf: x = 16'h2a0e; 12'h6c0: x = 16'h2a0a; 12'h6c1: x = 16'h2a07; 12'h6c2: x = 16'h2a03; 12'h6c3: x = 16'h29ff; 12'h6c4: x = 16'h29fc; 12'h6c5: x = 16'h29f8; 12'h6c6: x = 16'h29f5; 12'h6c7: x = 16'h29f1; 12'h6c8: x = 16'h29ed; 12'h6c9: x = 16'h29ea; 12'h6ca: x = 16'h29e6; 12'h6cb: x = 16'h29e3; 12'h6cc: x = 16'h29df; 12'h6cd: x = 16'h29db; 12'h6ce: x = 16'h29d8; 12'h6cf: x = 16'h29d4; 12'h6d0: x = 16'h29d1; 12'h6d1: x = 16'h29cd; 12'h6d2: x = 16'h29c9; 12'h6d3: x = 16'h29c6; 12'h6d4: x = 16'h29c2; 12'h6d5: x = 16'h29bf; 12'h6d6: x = 16'h29bb; 12'h6d7: x = 16'h29b7; 12'h6d8: x = 16'h29b4; 12'h6d9: x = 16'h29b0; 12'h6da: x = 16'h29ad; 12'h6db: x = 16'h29a9; 12'h6dc: x = 16'h29a6; 12'h6dd: x = 16'h29a2; 12'h6de: x = 16'h299e; 12'h6df: x = 16'h299b; 12'h6e0: x = 16'h2997; 12'h6e1: x = 16'h2994; 12'h6e2: x = 16'h2990; 12'h6e3: x = 16'h298c; 12'h6e4: x = 16'h2989; 12'h6e5: x = 16'h2985; 12'h6e6: x = 16'h2982; 12'h6e7: x = 16'h297e; 12'h6e8: x = 16'h297b; 12'h6e9: x = 16'h2977; 12'h6ea: x = 16'h2973; 12'h6eb: x = 16'h2970; 12'h6ec: x = 16'h296c; 12'h6ed: x = 16'h2969; 12'h6ee: x = 16'h2965; 12'h6ef: x = 16'h2962; 12'h6f0: x = 16'h295e; 12'h6f1: x = 16'h295a; 12'h6f2: x = 16'h2957; 12'h6f3: x = 16'h2953; 12'h6f4: x = 16'h2950; 12'h6f5: x = 16'h294c; 12'h6f6: x = 16'h2949; 12'h6f7: x = 16'h2945; 12'h6f8: x = 16'h2941; 12'h6f9: x = 16'h293e; 12'h6fa: x = 16'h293a; 12'h6fb: x = 16'h2937; 12'h6fc: x = 16'h2933; 12'h6fd: x = 16'h2930; 12'h6fe: x = 16'h292c; 12'h6ff: x = 16'h2929; 12'h700: x = 16'h2925; 12'h701: x = 16'h2921; 12'h702: x = 16'h291e; 12'h703: x = 16'h291a; 12'h704: x = 16'h2917; 12'h705: x = 16'h2913; 12'h706: x = 16'h2910; 12'h707: x = 16'h290c; 12'h708: x = 16'h2909; 12'h709: x = 16'h2905; 12'h70a: x = 16'h2902; 12'h70b: x = 16'h28fe; 12'h70c: x = 16'h28fa; 12'h70d: x = 16'h28f7; 12'h70e: x = 16'h28f3; 12'h70f: x = 16'h28f0; 12'h710: x = 16'h28ec; 12'h711: x = 16'h28e9; 12'h712: x = 16'h28e5; 12'h713: x = 16'h28e2; 12'h714: x = 16'h28de; 12'h715: x = 16'h28db; 12'h716: x = 16'h28d7; 12'h717: x = 16'h28d3; 12'h718: x = 16'h28d0; 12'h719: x = 16'h28cc; 12'h71a: x = 16'h28c9; 12'h71b: x = 16'h28c5; 12'h71c: x = 16'h28c2; 12'h71d: x = 16'h28be; 12'h71e: x = 16'h28bb; 12'h71f: x = 16'h28b7; 12'h720: x = 16'h28b4; 12'h721: x = 16'h28b0; 12'h722: x = 16'h28ad; 12'h723: x = 16'h28a9; 12'h724: x = 16'h28a6; 12'h725: x = 16'h28a2; 12'h726: x = 16'h289e; 12'h727: x = 16'h289b; 12'h728: x = 16'h2897; 12'h729: x = 16'h2894; 12'h72a: x = 16'h2890; 12'h72b: x = 16'h288d; 12'h72c: x = 16'h2889; 12'h72d: x = 16'h2886; 12'h72e: x = 16'h2882; 12'h72f: x = 16'h287f; 12'h730: x = 16'h287b; 12'h731: x = 16'h2878; 12'h732: x = 16'h2874; 12'h733: x = 16'h2871; 12'h734: x = 16'h286d; 12'h735: x = 16'h286a; 12'h736: x = 16'h2866; 12'h737: x = 16'h2863; 12'h738: x = 16'h285f; 12'h739: x = 16'h285c; 12'h73a: x = 16'h2858; 12'h73b: x = 16'h2855; 12'h73c: x = 16'h2851; 12'h73d: x = 16'h284e; 12'h73e: x = 16'h284a; 12'h73f: x = 16'h2847; 12'h740: x = 16'h2843; 12'h741: x = 16'h2840; 12'h742: x = 16'h283c; 12'h743: x = 16'h2839; 12'h744: x = 16'h2835; 12'h745: x = 16'h2831; 12'h746: x = 16'h282e; 12'h747: x = 16'h282a; 12'h748: x = 16'h2827; 12'h749: x = 16'h2823; 12'h74a: x = 16'h2820; 12'h74b: x = 16'h281c; 12'h74c: x = 16'h2819; 12'h74d: x = 16'h2815; 12'h74e: x = 16'h2812; 12'h74f: x = 16'h280e; 12'h750: x = 16'h280b; 12'h751: x = 16'h2807; 12'h752: x = 16'h2804; 12'h753: x = 16'h2800; 12'h754: x = 16'h27fd; 12'h755: x = 16'h27fa; 12'h756: x = 16'h27f6; 12'h757: x = 16'h27f3; 12'h758: x = 16'h27ef; 12'h759: x = 16'h27ec; 12'h75a: x = 16'h27e8; 12'h75b: x = 16'h27e5; 12'h75c: x = 16'h27e1; 12'h75d: x = 16'h27de; 12'h75e: x = 16'h27da; 12'h75f: x = 16'h27d7; 12'h760: x = 16'h27d3; 12'h761: x = 16'h27d0; 12'h762: x = 16'h27cc; 12'h763: x = 16'h27c9; 12'h764: x = 16'h27c5; 12'h765: x = 16'h27c2; 12'h766: x = 16'h27be; 12'h767: x = 16'h27bb; 12'h768: x = 16'h27b7; 12'h769: x = 16'h27b4; 12'h76a: x = 16'h27b0; 12'h76b: x = 16'h27ad; 12'h76c: x = 16'h27a9; 12'h76d: x = 16'h27a6; 12'h76e: x = 16'h27a2; 12'h76f: x = 16'h279f; 12'h770: x = 16'h279b; 12'h771: x = 16'h2798; 12'h772: x = 16'h2794; 12'h773: x = 16'h2791; 12'h774: x = 16'h278e; 12'h775: x = 16'h278a; 12'h776: x = 16'h2787; 12'h777: x = 16'h2783; 12'h778: x = 16'h2780; 12'h779: x = 16'h277c; 12'h77a: x = 16'h2779; 12'h77b: x = 16'h2775; 12'h77c: x = 16'h2772; 12'h77d: x = 16'h276e; 12'h77e: x = 16'h276b; 12'h77f: x = 16'h2767; 12'h780: x = 16'h2764; 12'h781: x = 16'h2760; 12'h782: x = 16'h275d; 12'h783: x = 16'h2759; 12'h784: x = 16'h2756; 12'h785: x = 16'h2753; 12'h786: x = 16'h274f; 12'h787: x = 16'h274c; 12'h788: x = 16'h2748; 12'h789: x = 16'h2745; 12'h78a: x = 16'h2741; 12'h78b: x = 16'h273e; 12'h78c: x = 16'h273a; 12'h78d: x = 16'h2737; 12'h78e: x = 16'h2733; 12'h78f: x = 16'h2730; 12'h790: x = 16'h272d; 12'h791: x = 16'h2729; 12'h792: x = 16'h2726; 12'h793: x = 16'h2722; 12'h794: x = 16'h271f; 12'h795: x = 16'h271b; 12'h796: x = 16'h2718; 12'h797: x = 16'h2714; 12'h798: x = 16'h2711; 12'h799: x = 16'h270d; 12'h79a: x = 16'h270a; 12'h79b: x = 16'h2707; 12'h79c: x = 16'h2703; 12'h79d: x = 16'h2700; 12'h79e: x = 16'h26fc; 12'h79f: x = 16'h26f9; 12'h7a0: x = 16'h26f5; 12'h7a1: x = 16'h26f2; 12'h7a2: x = 16'h26ee; 12'h7a3: x = 16'h26eb; 12'h7a4: x = 16'h26e7; 12'h7a5: x = 16'h26e4; 12'h7a6: x = 16'h26e1; 12'h7a7: x = 16'h26dd; 12'h7a8: x = 16'h26da; 12'h7a9: x = 16'h26d6; 12'h7aa: x = 16'h26d3; 12'h7ab: x = 16'h26cf; 12'h7ac: x = 16'h26cc; 12'h7ad: x = 16'h26c9; 12'h7ae: x = 16'h26c5; 12'h7af: x = 16'h26c2; 12'h7b0: x = 16'h26be; 12'h7b1: x = 16'h26bb; 12'h7b2: x = 16'h26b7; 12'h7b3: x = 16'h26b4; 12'h7b4: x = 16'h26b0; 12'h7b5: x = 16'h26ad; 12'h7b6: x = 16'h26aa; 12'h7b7: x = 16'h26a6; 12'h7b8: x = 16'h26a3; 12'h7b9: x = 16'h269f; 12'h7ba: x = 16'h269c; 12'h7bb: x = 16'h2698; 12'h7bc: x = 16'h2695; 12'h7bd: x = 16'h2692; 12'h7be: x = 16'h268e; 12'h7bf: x = 16'h268b; 12'h7c0: x = 16'h2687; 12'h7c1: x = 16'h2684; 12'h7c2: x = 16'h2680; 12'h7c3: x = 16'h267d; 12'h7c4: x = 16'h267a; 12'h7c5: x = 16'h2676; 12'h7c6: x = 16'h2673; 12'h7c7: x = 16'h266f; 12'h7c8: x = 16'h266c; 12'h7c9: x = 16'h2668; 12'h7ca: x = 16'h2665; 12'h7cb: x = 16'h2662; 12'h7cc: x = 16'h265e; 12'h7cd: x = 16'h265b; 12'h7ce: x = 16'h2657; 12'h7cf: x = 16'h2654; 12'h7d0: x = 16'h2650; 12'h7d1: x = 16'h264d; 12'h7d2: x = 16'h264a; 12'h7d3: x = 16'h2646; 12'h7d4: x = 16'h2643; 12'h7d5: x = 16'h263f; 12'h7d6: x = 16'h263c; 12'h7d7: x = 16'h2639; 12'h7d8: x = 16'h2635; 12'h7d9: x = 16'h2632; 12'h7da: x = 16'h262e; 12'h7db: x = 16'h262b; 12'h7dc: x = 16'h2627; 12'h7dd: x = 16'h2624; 12'h7de: x = 16'h2621; 12'h7df: x = 16'h261d; 12'h7e0: x = 16'h261a; 12'h7e1: x = 16'h2616; 12'h7e2: x = 16'h2613; 12'h7e3: x = 16'h2610; 12'h7e4: x = 16'h260c; 12'h7e5: x = 16'h2609; 12'h7e6: x = 16'h2605; 12'h7e7: x = 16'h2602; 12'h7e8: x = 16'h25ff; 12'h7e9: x = 16'h25fb; 12'h7ea: x = 16'h25f8; 12'h7eb: x = 16'h25f4; 12'h7ec: x = 16'h25f1; 12'h7ed: x = 16'h25ed; 12'h7ee: x = 16'h25ea; 12'h7ef: x = 16'h25e7; 12'h7f0: x = 16'h25e3; 12'h7f1: x = 16'h25e0; 12'h7f2: x = 16'h25dc; 12'h7f3: x = 16'h25d9; 12'h7f4: x = 16'h25d6; 12'h7f5: x = 16'h25d2; 12'h7f6: x = 16'h25cf; 12'h7f7: x = 16'h25cb; 12'h7f8: x = 16'h25c8; 12'h7f9: x = 16'h25c5; 12'h7fa: x = 16'h25c1; 12'h7fb: x = 16'h25be; 12'h7fc: x = 16'h25ba; 12'h7fd: x = 16'h25b7; 12'h7fe: x = 16'h25b4; 12'h7ff: x = 16'h25b0; 12'h800: x = 16'h25ad; 12'h801: x = 16'h25a9; 12'h802: x = 16'h25a6; 12'h803: x = 16'h25a3; 12'h804: x = 16'h259f; 12'h805: x = 16'h259c; 12'h806: x = 16'h2598; 12'h807: x = 16'h2595; 12'h808: x = 16'h2592; 12'h809: x = 16'h258e; 12'h80a: x = 16'h258b; 12'h80b: x = 16'h2588; 12'h80c: x = 16'h2584; 12'h80d: x = 16'h2581; 12'h80e: x = 16'h257d; 12'h80f: x = 16'h257a; 12'h810: x = 16'h2577; 12'h811: x = 16'h2573; 12'h812: x = 16'h2570; 12'h813: x = 16'h256c; 12'h814: x = 16'h2569; 12'h815: x = 16'h2566; 12'h816: x = 16'h2562; 12'h817: x = 16'h255f; 12'h818: x = 16'h255b; 12'h819: x = 16'h2558; 12'h81a: x = 16'h2555; 12'h81b: x = 16'h2551; 12'h81c: x = 16'h254e; 12'h81d: x = 16'h254b; 12'h81e: x = 16'h2547; 12'h81f: x = 16'h2544; 12'h820: x = 16'h2540; 12'h821: x = 16'h253d; 12'h822: x = 16'h253a; 12'h823: x = 16'h2536; 12'h824: x = 16'h2533; 12'h825: x = 16'h252f; 12'h826: x = 16'h252c; 12'h827: x = 16'h2529; 12'h828: x = 16'h2525; 12'h829: x = 16'h2522; 12'h82a: x = 16'h251f; 12'h82b: x = 16'h251b; 12'h82c: x = 16'h2518; 12'h82d: x = 16'h2514; 12'h82e: x = 16'h2511; 12'h82f: x = 16'h250e; 12'h830: x = 16'h250a; 12'h831: x = 16'h2507; 12'h832: x = 16'h2504; 12'h833: x = 16'h2500; 12'h834: x = 16'h24fd; 12'h835: x = 16'h24f9; 12'h836: x = 16'h24f6; 12'h837: x = 16'h24f3; 12'h838: x = 16'h24ef; 12'h839: x = 16'h24ec; 12'h83a: x = 16'h24e9; 12'h83b: x = 16'h24e5; 12'h83c: x = 16'h24e2; 12'h83d: x = 16'h24de; 12'h83e: x = 16'h24db; 12'h83f: x = 16'h24d8; 12'h840: x = 16'h24d4; 12'h841: x = 16'h24d1; 12'h842: x = 16'h24ce; 12'h843: x = 16'h24ca; 12'h844: x = 16'h24c7; 12'h845: x = 16'h24c3; 12'h846: x = 16'h24c0; 12'h847: x = 16'h24bd; 12'h848: x = 16'h24b9; 12'h849: x = 16'h24b6; 12'h84a: x = 16'h24b3; 12'h84b: x = 16'h24af; 12'h84c: x = 16'h24ac; 12'h84d: x = 16'h24a9; 12'h84e: x = 16'h24a5; 12'h84f: x = 16'h24a2; 12'h850: x = 16'h249e; 12'h851: x = 16'h249b; 12'h852: x = 16'h2498; 12'h853: x = 16'h2494; 12'h854: x = 16'h2491; 12'h855: x = 16'h248e; 12'h856: x = 16'h248a; 12'h857: x = 16'h2487; 12'h858: x = 16'h2484; 12'h859: x = 16'h2480; 12'h85a: x = 16'h247d; 12'h85b: x = 16'h2479; 12'h85c: x = 16'h2476; 12'h85d: x = 16'h2473; 12'h85e: x = 16'h246f; 12'h85f: x = 16'h246c; 12'h860: x = 16'h2469; 12'h861: x = 16'h2465; 12'h862: x = 16'h2462; 12'h863: x = 16'h245f; 12'h864: x = 16'h245b; 12'h865: x = 16'h2458; 12'h866: x = 16'h2455; 12'h867: x = 16'h2451; 12'h868: x = 16'h244e; 12'h869: x = 16'h244a; 12'h86a: x = 16'h2447; 12'h86b: x = 16'h2444; 12'h86c: x = 16'h2440; 12'h86d: x = 16'h243d; 12'h86e: x = 16'h243a; 12'h86f: x = 16'h2436; 12'h870: x = 16'h2433; 12'h871: x = 16'h2430; 12'h872: x = 16'h242c; 12'h873: x = 16'h2429; 12'h874: x = 16'h2426; 12'h875: x = 16'h2422; 12'h876: x = 16'h241f; 12'h877: x = 16'h241c; 12'h878: x = 16'h2418; 12'h879: x = 16'h2415; 12'h87a: x = 16'h2411; 12'h87b: x = 16'h240e; 12'h87c: x = 16'h240b; 12'h87d: x = 16'h2407; 12'h87e: x = 16'h2404; 12'h87f: x = 16'h2401; 12'h880: x = 16'h23fd; 12'h881: x = 16'h23fa; 12'h882: x = 16'h23f7; 12'h883: x = 16'h23f3; 12'h884: x = 16'h23f0; 12'h885: x = 16'h23ed; 12'h886: x = 16'h23e9; 12'h887: x = 16'h23e6; 12'h888: x = 16'h23e3; 12'h889: x = 16'h23df; 12'h88a: x = 16'h23dc; 12'h88b: x = 16'h23d9; 12'h88c: x = 16'h23d5; 12'h88d: x = 16'h23d2; 12'h88e: x = 16'h23cf; 12'h88f: x = 16'h23cb; 12'h890: x = 16'h23c8; 12'h891: x = 16'h23c5; 12'h892: x = 16'h23c1; 12'h893: x = 16'h23be; 12'h894: x = 16'h23bb; 12'h895: x = 16'h23b7; 12'h896: x = 16'h23b4; 12'h897: x = 16'h23b0; 12'h898: x = 16'h23ad; 12'h899: x = 16'h23aa; 12'h89a: x = 16'h23a6; 12'h89b: x = 16'h23a3; 12'h89c: x = 16'h23a0; 12'h89d: x = 16'h239c; 12'h89e: x = 16'h2399; 12'h89f: x = 16'h2396; 12'h8a0: x = 16'h2392; 12'h8a1: x = 16'h238f; 12'h8a2: x = 16'h238c; 12'h8a3: x = 16'h2388; 12'h8a4: x = 16'h2385; 12'h8a5: x = 16'h2382; 12'h8a6: x = 16'h237e; 12'h8a7: x = 16'h237b; 12'h8a8: x = 16'h2378; 12'h8a9: x = 16'h2374; 12'h8aa: x = 16'h2371; 12'h8ab: x = 16'h236e; 12'h8ac: x = 16'h236a; 12'h8ad: x = 16'h2367; 12'h8ae: x = 16'h2364; 12'h8af: x = 16'h2360; 12'h8b0: x = 16'h235d; 12'h8b1: x = 16'h235a; 12'h8b2: x = 16'h2356; 12'h8b3: x = 16'h2353; 12'h8b4: x = 16'h2350; 12'h8b5: x = 16'h234c; 12'h8b6: x = 16'h2349; 12'h8b7: x = 16'h2346; 12'h8b8: x = 16'h2342; 12'h8b9: x = 16'h233f; 12'h8ba: x = 16'h233c; 12'h8bb: x = 16'h2338; 12'h8bc: x = 16'h2335; 12'h8bd: x = 16'h2332; 12'h8be: x = 16'h232e; 12'h8bf: x = 16'h232b; 12'h8c0: x = 16'h2328; 12'h8c1: x = 16'h2324; 12'h8c2: x = 16'h2321; 12'h8c3: x = 16'h231e; 12'h8c4: x = 16'h231a; 12'h8c5: x = 16'h2317; 12'h8c6: x = 16'h2314; 12'h8c7: x = 16'h2310; 12'h8c8: x = 16'h230d; 12'h8c9: x = 16'h230a; 12'h8ca: x = 16'h2307; 12'h8cb: x = 16'h2303; 12'h8cc: x = 16'h2300; 12'h8cd: x = 16'h22fd; 12'h8ce: x = 16'h22f9; 12'h8cf: x = 16'h22f6; 12'h8d0: x = 16'h22f3; 12'h8d1: x = 16'h22ef; 12'h8d2: x = 16'h22ec; 12'h8d3: x = 16'h22e9; 12'h8d4: x = 16'h22e5; 12'h8d5: x = 16'h22e2; 12'h8d6: x = 16'h22df; 12'h8d7: x = 16'h22db; 12'h8d8: x = 16'h22d8; 12'h8d9: x = 16'h22d5; 12'h8da: x = 16'h22d1; 12'h8db: x = 16'h22ce; 12'h8dc: x = 16'h22cb; 12'h8dd: x = 16'h22c7; 12'h8de: x = 16'h22c4; 12'h8df: x = 16'h22c1; 12'h8e0: x = 16'h22bd; 12'h8e1: x = 16'h22ba; 12'h8e2: x = 16'h22b7; 12'h8e3: x = 16'h22b3; 12'h8e4: x = 16'h22b0; 12'h8e5: x = 16'h22ad; 12'h8e6: x = 16'h22a9; 12'h8e7: x = 16'h22a6; 12'h8e8: x = 16'h22a3; 12'h8e9: x = 16'h22a0; 12'h8ea: x = 16'h229c; 12'h8eb: x = 16'h2299; 12'h8ec: x = 16'h2296; 12'h8ed: x = 16'h2292; 12'h8ee: x = 16'h228f; 12'h8ef: x = 16'h228c; 12'h8f0: x = 16'h2288; 12'h8f1: x = 16'h2285; 12'h8f2: x = 16'h2282; 12'h8f3: x = 16'h227e; 12'h8f4: x = 16'h227b; 12'h8f5: x = 16'h2278; 12'h8f6: x = 16'h2274; 12'h8f7: x = 16'h2271; 12'h8f8: x = 16'h226e; 12'h8f9: x = 16'h226a; 12'h8fa: x = 16'h2267; 12'h8fb: x = 16'h2264; 12'h8fc: x = 16'h2260; 12'h8fd: x = 16'h225d; 12'h8fe: x = 16'h225a; 12'h8ff: x = 16'h2257; 12'h900: x = 16'h2253; 12'h901: x = 16'h2250; 12'h902: x = 16'h224d; 12'h903: x = 16'h2249; 12'h904: x = 16'h2246; 12'h905: x = 16'h2243; 12'h906: x = 16'h223f; 12'h907: x = 16'h223c; 12'h908: x = 16'h2239; 12'h909: x = 16'h2235; 12'h90a: x = 16'h2232; 12'h90b: x = 16'h222f; 12'h90c: x = 16'h222b; 12'h90d: x = 16'h2228; 12'h90e: x = 16'h2225; 12'h90f: x = 16'h2222; 12'h910: x = 16'h221e; 12'h911: x = 16'h221b; 12'h912: x = 16'h2218; 12'h913: x = 16'h2214; 12'h914: x = 16'h2211; 12'h915: x = 16'h220e; 12'h916: x = 16'h220a; 12'h917: x = 16'h2207; 12'h918: x = 16'h2204; 12'h919: x = 16'h2200; 12'h91a: x = 16'h21fd; 12'h91b: x = 16'h21fa; 12'h91c: x = 16'h21f6; 12'h91d: x = 16'h21f3; 12'h91e: x = 16'h21f0; 12'h91f: x = 16'h21ed; 12'h920: x = 16'h21e9; 12'h921: x = 16'h21e6; 12'h922: x = 16'h21e3; 12'h923: x = 16'h21df; 12'h924: x = 16'h21dc; 12'h925: x = 16'h21d9; 12'h926: x = 16'h21d5; 12'h927: x = 16'h21d2; 12'h928: x = 16'h21cf; 12'h929: x = 16'h21cb; 12'h92a: x = 16'h21c8; 12'h92b: x = 16'h21c5; 12'h92c: x = 16'h21c2; 12'h92d: x = 16'h21be; 12'h92e: x = 16'h21bb; 12'h92f: x = 16'h21b8; 12'h930: x = 16'h21b4; 12'h931: x = 16'h21b1; 12'h932: x = 16'h21ae; 12'h933: x = 16'h21aa; 12'h934: x = 16'h21a7; 12'h935: x = 16'h21a4; 12'h936: x = 16'h21a0; 12'h937: x = 16'h219d; 12'h938: x = 16'h219a; 12'h939: x = 16'h2197; 12'h93a: x = 16'h2193; 12'h93b: x = 16'h2190; 12'h93c: x = 16'h218d; 12'h93d: x = 16'h2189; 12'h93e: x = 16'h2186; 12'h93f: x = 16'h2183; 12'h940: x = 16'h217f; 12'h941: x = 16'h217c; 12'h942: x = 16'h2179; 12'h943: x = 16'h2176; 12'h944: x = 16'h2172; 12'h945: x = 16'h216f; 12'h946: x = 16'h216c; 12'h947: x = 16'h2168; 12'h948: x = 16'h2165; 12'h949: x = 16'h2162; 12'h94a: x = 16'h215e; 12'h94b: x = 16'h215b; 12'h94c: x = 16'h2158; 12'h94d: x = 16'h2154; 12'h94e: x = 16'h2151; 12'h94f: x = 16'h214e; 12'h950: x = 16'h214b; 12'h951: x = 16'h2147; 12'h952: x = 16'h2144; 12'h953: x = 16'h2141; 12'h954: x = 16'h213d; 12'h955: x = 16'h213a; 12'h956: x = 16'h2137; 12'h957: x = 16'h2133; 12'h958: x = 16'h2130; 12'h959: x = 16'h212d; 12'h95a: x = 16'h212a; 12'h95b: x = 16'h2126; 12'h95c: x = 16'h2123; 12'h95d: x = 16'h2120; 12'h95e: x = 16'h211c; 12'h95f: x = 16'h2119; 12'h960: x = 16'h2116; 12'h961: x = 16'h2112; 12'h962: x = 16'h210f; 12'h963: x = 16'h210c; 12'h964: x = 16'h2109; 12'h965: x = 16'h2105; 12'h966: x = 16'h2102; 12'h967: x = 16'h20ff; 12'h968: x = 16'h20fb; 12'h969: x = 16'h20f8; 12'h96a: x = 16'h20f5; 12'h96b: x = 16'h20f1; 12'h96c: x = 16'h20ee; 12'h96d: x = 16'h20eb; 12'h96e: x = 16'h20e8; 12'h96f: x = 16'h20e4; 12'h970: x = 16'h20e1; 12'h971: x = 16'h20de; 12'h972: x = 16'h20da; 12'h973: x = 16'h20d7; 12'h974: x = 16'h20d4; 12'h975: x = 16'h20d0; 12'h976: x = 16'h20cd; 12'h977: x = 16'h20ca; 12'h978: x = 16'h20c7; 12'h979: x = 16'h20c3; 12'h97a: x = 16'h20c0; 12'h97b: x = 16'h20bd; 12'h97c: x = 16'h20b9; 12'h97d: x = 16'h20b6; 12'h97e: x = 16'h20b3; 12'h97f: x = 16'h20af; 12'h980: x = 16'h20ac; 12'h981: x = 16'h20a9; 12'h982: x = 16'h20a6; 12'h983: x = 16'h20a2; 12'h984: x = 16'h209f; 12'h985: x = 16'h209c; 12'h986: x = 16'h2098; 12'h987: x = 16'h2095; 12'h988: x = 16'h2092; 12'h989: x = 16'h208e; 12'h98a: x = 16'h208b; 12'h98b: x = 16'h2088; 12'h98c: x = 16'h2085; 12'h98d: x = 16'h2081; 12'h98e: x = 16'h207e; 12'h98f: x = 16'h207b; 12'h990: x = 16'h2077; 12'h991: x = 16'h2074; 12'h992: x = 16'h2071; 12'h993: x = 16'h206d; 12'h994: x = 16'h206a; 12'h995: x = 16'h2067; 12'h996: x = 16'h2064; 12'h997: x = 16'h2060; 12'h998: x = 16'h205d; 12'h999: x = 16'h205a; 12'h99a: x = 16'h2056; 12'h99b: x = 16'h2053; 12'h99c: x = 16'h2050; 12'h99d: x = 16'h204c; 12'h99e: x = 16'h2049; 12'h99f: x = 16'h2046; 12'h9a0: x = 16'h2043; 12'h9a1: x = 16'h203f; 12'h9a2: x = 16'h203c; 12'h9a3: x = 16'h2039; 12'h9a4: x = 16'h2035; 12'h9a5: x = 16'h2032; 12'h9a6: x = 16'h202f; 12'h9a7: x = 16'h202c; 12'h9a8: x = 16'h2028; 12'h9a9: x = 16'h2025; 12'h9aa: x = 16'h2022; 12'h9ab: x = 16'h201e; 12'h9ac: x = 16'h201b; 12'h9ad: x = 16'h2018; 12'h9ae: x = 16'h2014; 12'h9af: x = 16'h2011; 12'h9b0: x = 16'h200e; 12'h9b1: x = 16'h200b; 12'h9b2: x = 16'h2007; 12'h9b3: x = 16'h2004; 12'h9b4: x = 16'h2001; 12'h9b5: x = 16'h1ffd; 12'h9b6: x = 16'h1ffa; 12'h9b7: x = 16'h1ff7; 12'h9b8: x = 16'h1ff3; 12'h9b9: x = 16'h1ff0; 12'h9ba: x = 16'h1fed; 12'h9bb: x = 16'h1fea; 12'h9bc: x = 16'h1fe6; 12'h9bd: x = 16'h1fe3; 12'h9be: x = 16'h1fe0; 12'h9bf: x = 16'h1fdc; 12'h9c0: x = 16'h1fd9; 12'h9c1: x = 16'h1fd6; 12'h9c2: x = 16'h1fd2; 12'h9c3: x = 16'h1fcf; 12'h9c4: x = 16'h1fcc; 12'h9c5: x = 16'h1fc9; 12'h9c6: x = 16'h1fc5; 12'h9c7: x = 16'h1fc2; 12'h9c8: x = 16'h1fbf; 12'h9c9: x = 16'h1fbb; 12'h9ca: x = 16'h1fb8; 12'h9cb: x = 16'h1fb5; 12'h9cc: x = 16'h1fb2; 12'h9cd: x = 16'h1fae; 12'h9ce: x = 16'h1fab; 12'h9cf: x = 16'h1fa8; 12'h9d0: x = 16'h1fa4; 12'h9d1: x = 16'h1fa1; 12'h9d2: x = 16'h1f9e; 12'h9d3: x = 16'h1f9a; 12'h9d4: x = 16'h1f97; 12'h9d5: x = 16'h1f94; 12'h9d6: x = 16'h1f91; 12'h9d7: x = 16'h1f8d; 12'h9d8: x = 16'h1f8a; 12'h9d9: x = 16'h1f87; 12'h9da: x = 16'h1f83; 12'h9db: x = 16'h1f80; 12'h9dc: x = 16'h1f7d; 12'h9dd: x = 16'h1f79; 12'h9de: x = 16'h1f76; 12'h9df: x = 16'h1f73; 12'h9e0: x = 16'h1f70; 12'h9e1: x = 16'h1f6c; 12'h9e2: x = 16'h1f69; 12'h9e3: x = 16'h1f66; 12'h9e4: x = 16'h1f62; 12'h9e5: x = 16'h1f5f; 12'h9e6: x = 16'h1f5c; 12'h9e7: x = 16'h1f58; 12'h9e8: x = 16'h1f55; 12'h9e9: x = 16'h1f52; 12'h9ea: x = 16'h1f4f; 12'h9eb: x = 16'h1f4b; 12'h9ec: x = 16'h1f48; 12'h9ed: x = 16'h1f45; 12'h9ee: x = 16'h1f41; 12'h9ef: x = 16'h1f3e; 12'h9f0: x = 16'h1f3b; 12'h9f1: x = 16'h1f37; 12'h9f2: x = 16'h1f34; 12'h9f3: x = 16'h1f31; 12'h9f4: x = 16'h1f2e; 12'h9f5: x = 16'h1f2a; 12'h9f6: x = 16'h1f27; 12'h9f7: x = 16'h1f24; 12'h9f8: x = 16'h1f20; 12'h9f9: x = 16'h1f1d; 12'h9fa: x = 16'h1f1a; 12'h9fb: x = 16'h1f16; 12'h9fc: x = 16'h1f13; 12'h9fd: x = 16'h1f10; 12'h9fe: x = 16'h1f0d; 12'h9ff: x = 16'h1f09; 12'ha00: x = 16'h1f06; 12'ha01: x = 16'h1f03; 12'ha02: x = 16'h1eff; 12'ha03: x = 16'h1efc; 12'ha04: x = 16'h1ef9; 12'ha05: x = 16'h1ef5; 12'ha06: x = 16'h1ef2; 12'ha07: x = 16'h1eef; 12'ha08: x = 16'h1eec; 12'ha09: x = 16'h1ee8; 12'ha0a: x = 16'h1ee5; 12'ha0b: x = 16'h1ee2; 12'ha0c: x = 16'h1ede; 12'ha0d: x = 16'h1edb; 12'ha0e: x = 16'h1ed8; 12'ha0f: x = 16'h1ed4; 12'ha10: x = 16'h1ed1; 12'ha11: x = 16'h1ece; 12'ha12: x = 16'h1ecb; 12'ha13: x = 16'h1ec7; 12'ha14: x = 16'h1ec4; 12'ha15: x = 16'h1ec1; 12'ha16: x = 16'h1ebd; 12'ha17: x = 16'h1eba; 12'ha18: x = 16'h1eb7; 12'ha19: x = 16'h1eb3; 12'ha1a: x = 16'h1eb0; 12'ha1b: x = 16'h1ead; 12'ha1c: x = 16'h1eaa; 12'ha1d: x = 16'h1ea6; 12'ha1e: x = 16'h1ea3; 12'ha1f: x = 16'h1ea0; 12'ha20: x = 16'h1e9c; 12'ha21: x = 16'h1e99; 12'ha22: x = 16'h1e96; 12'ha23: x = 16'h1e92; 12'ha24: x = 16'h1e8f; 12'ha25: x = 16'h1e8c; 12'ha26: x = 16'h1e88; 12'ha27: x = 16'h1e85; 12'ha28: x = 16'h1e82; 12'ha29: x = 16'h1e7f; 12'ha2a: x = 16'h1e7b; 12'ha2b: x = 16'h1e78; 12'ha2c: x = 16'h1e75; 12'ha2d: x = 16'h1e71; 12'ha2e: x = 16'h1e6e; 12'ha2f: x = 16'h1e6b; 12'ha30: x = 16'h1e67; 12'ha31: x = 16'h1e64; 12'ha32: x = 16'h1e61; 12'ha33: x = 16'h1e5e; 12'ha34: x = 16'h1e5a; 12'ha35: x = 16'h1e57; 12'ha36: x = 16'h1e54; 12'ha37: x = 16'h1e50; 12'ha38: x = 16'h1e4d; 12'ha39: x = 16'h1e4a; 12'ha3a: x = 16'h1e46; 12'ha3b: x = 16'h1e43; 12'ha3c: x = 16'h1e40; 12'ha3d: x = 16'h1e3c; 12'ha3e: x = 16'h1e39; 12'ha3f: x = 16'h1e36; 12'ha40: x = 16'h1e33; 12'ha41: x = 16'h1e2f; 12'ha42: x = 16'h1e2c; 12'ha43: x = 16'h1e29; 12'ha44: x = 16'h1e25; 12'ha45: x = 16'h1e22; 12'ha46: x = 16'h1e1f; 12'ha47: x = 16'h1e1b; 12'ha48: x = 16'h1e18; 12'ha49: x = 16'h1e15; 12'ha4a: x = 16'h1e11; 12'ha4b: x = 16'h1e0e; 12'ha4c: x = 16'h1e0b; 12'ha4d: x = 16'h1e07; 12'ha4e: x = 16'h1e04; 12'ha4f: x = 16'h1e01; 12'ha50: x = 16'h1dfe; 12'ha51: x = 16'h1dfa; 12'ha52: x = 16'h1df7; 12'ha53: x = 16'h1df4; 12'ha54: x = 16'h1df0; 12'ha55: x = 16'h1ded; 12'ha56: x = 16'h1dea; 12'ha57: x = 16'h1de6; 12'ha58: x = 16'h1de3; 12'ha59: x = 16'h1de0; 12'ha5a: x = 16'h1ddc; 12'ha5b: x = 16'h1dd9; 12'ha5c: x = 16'h1dd6; 12'ha5d: x = 16'h1dd3; 12'ha5e: x = 16'h1dcf; 12'ha5f: x = 16'h1dcc; 12'ha60: x = 16'h1dc9; 12'ha61: x = 16'h1dc5; 12'ha62: x = 16'h1dc2; 12'ha63: x = 16'h1dbf; 12'ha64: x = 16'h1dbb; 12'ha65: x = 16'h1db8; 12'ha66: x = 16'h1db5; 12'ha67: x = 16'h1db1; 12'ha68: x = 16'h1dae; 12'ha69: x = 16'h1dab; 12'ha6a: x = 16'h1da7; 12'ha6b: x = 16'h1da4; 12'ha6c: x = 16'h1da1; 12'ha6d: x = 16'h1d9d; 12'ha6e: x = 16'h1d9a; 12'ha6f: x = 16'h1d97; 12'ha70: x = 16'h1d94; 12'ha71: x = 16'h1d90; 12'ha72: x = 16'h1d8d; 12'ha73: x = 16'h1d8a; 12'ha74: x = 16'h1d86; 12'ha75: x = 16'h1d83; 12'ha76: x = 16'h1d80; 12'ha77: x = 16'h1d7c; 12'ha78: x = 16'h1d79; 12'ha79: x = 16'h1d76; 12'ha7a: x = 16'h1d72; 12'ha7b: x = 16'h1d6f; 12'ha7c: x = 16'h1d6c; 12'ha7d: x = 16'h1d68; 12'ha7e: x = 16'h1d65; 12'ha7f: x = 16'h1d62; 12'ha80: x = 16'h1d5e; 12'ha81: x = 16'h1d5b; 12'ha82: x = 16'h1d58; 12'ha83: x = 16'h1d54; 12'ha84: x = 16'h1d51; 12'ha85: x = 16'h1d4e; 12'ha86: x = 16'h1d4b; 12'ha87: x = 16'h1d47; 12'ha88: x = 16'h1d44; 12'ha89: x = 16'h1d41; 12'ha8a: x = 16'h1d3d; 12'ha8b: x = 16'h1d3a; 12'ha8c: x = 16'h1d37; 12'ha8d: x = 16'h1d33; 12'ha8e: x = 16'h1d30; 12'ha8f: x = 16'h1d2d; 12'ha90: x = 16'h1d29; 12'ha91: x = 16'h1d26; 12'ha92: x = 16'h1d23; 12'ha93: x = 16'h1d1f; 12'ha94: x = 16'h1d1c; 12'ha95: x = 16'h1d19; 12'ha96: x = 16'h1d15; 12'ha97: x = 16'h1d12; 12'ha98: x = 16'h1d0f; 12'ha99: x = 16'h1d0b; 12'ha9a: x = 16'h1d08; 12'ha9b: x = 16'h1d05; 12'ha9c: x = 16'h1d01; 12'ha9d: x = 16'h1cfe; 12'ha9e: x = 16'h1cfb; 12'ha9f: x = 16'h1cf7; 12'haa0: x = 16'h1cf4; 12'haa1: x = 16'h1cf1; 12'haa2: x = 16'h1ced; 12'haa3: x = 16'h1cea; 12'haa4: x = 16'h1ce7; 12'haa5: x = 16'h1ce3; 12'haa6: x = 16'h1ce0; 12'haa7: x = 16'h1cdd; 12'haa8: x = 16'h1cd9; 12'haa9: x = 16'h1cd6; 12'haaa: x = 16'h1cd3; 12'haab: x = 16'h1ccf; 12'haac: x = 16'h1ccc; 12'haad: x = 16'h1cc9; 12'haae: x = 16'h1cc5; 12'haaf: x = 16'h1cc2; 12'hab0: x = 16'h1cbf; 12'hab1: x = 16'h1cbb; 12'hab2: x = 16'h1cb8; 12'hab3: x = 16'h1cb5; 12'hab4: x = 16'h1cb1; 12'hab5: x = 16'h1cae; 12'hab6: x = 16'h1cab; 12'hab7: x = 16'h1ca7; 12'hab8: x = 16'h1ca4; 12'hab9: x = 16'h1ca1; 12'haba: x = 16'h1c9d; 12'habb: x = 16'h1c9a; 12'habc: x = 16'h1c97; 12'habd: x = 16'h1c93; 12'habe: x = 16'h1c90; 12'habf: x = 16'h1c8d; 12'hac0: x = 16'h1c89; 12'hac1: x = 16'h1c86; 12'hac2: x = 16'h1c83; 12'hac3: x = 16'h1c7f; 12'hac4: x = 16'h1c7c; 12'hac5: x = 16'h1c79; 12'hac6: x = 16'h1c75; 12'hac7: x = 16'h1c72; 12'hac8: x = 16'h1c6f; 12'hac9: x = 16'h1c6b; 12'haca: x = 16'h1c68; 12'hacb: x = 16'h1c65; 12'hacc: x = 16'h1c61; 12'hacd: x = 16'h1c5e; 12'hace: x = 16'h1c5b; 12'hacf: x = 16'h1c57; 12'had0: x = 16'h1c54; 12'had1: x = 16'h1c51; 12'had2: x = 16'h1c4d; 12'had3: x = 16'h1c4a; 12'had4: x = 16'h1c47; 12'had5: x = 16'h1c43; 12'had6: x = 16'h1c40; 12'had7: x = 16'h1c3d; 12'had8: x = 16'h1c39; 12'had9: x = 16'h1c36; 12'hada: x = 16'h1c33; 12'hadb: x = 16'h1c2f; 12'hadc: x = 16'h1c2c; 12'hadd: x = 16'h1c28; 12'hade: x = 16'h1c25; 12'hadf: x = 16'h1c22; 12'hae0: x = 16'h1c1e; 12'hae1: x = 16'h1c1b; 12'hae2: x = 16'h1c18; 12'hae3: x = 16'h1c14; 12'hae4: x = 16'h1c11; 12'hae5: x = 16'h1c0e; 12'hae6: x = 16'h1c0a; 12'hae7: x = 16'h1c07; 12'hae8: x = 16'h1c04; 12'hae9: x = 16'h1c00; 12'haea: x = 16'h1bfd; 12'haeb: x = 16'h1bfa; 12'haec: x = 16'h1bf6; 12'haed: x = 16'h1bf3; 12'haee: x = 16'h1bf0; 12'haef: x = 16'h1bec; 12'haf0: x = 16'h1be9; 12'haf1: x = 16'h1be5; 12'haf2: x = 16'h1be2; 12'haf3: x = 16'h1bdf; 12'haf4: x = 16'h1bdb; 12'haf5: x = 16'h1bd8; 12'haf6: x = 16'h1bd5; 12'haf7: x = 16'h1bd1; 12'haf8: x = 16'h1bce; 12'haf9: x = 16'h1bcb; 12'hafa: x = 16'h1bc7; 12'hafb: x = 16'h1bc4; 12'hafc: x = 16'h1bc1; 12'hafd: x = 16'h1bbd; 12'hafe: x = 16'h1bba; 12'haff: x = 16'h1bb6; 12'hb00: x = 16'h1bb3; 12'hb01: x = 16'h1bb0; 12'hb02: x = 16'h1bac; 12'hb03: x = 16'h1ba9; 12'hb04: x = 16'h1ba6; 12'hb05: x = 16'h1ba2; 12'hb06: x = 16'h1b9f; 12'hb07: x = 16'h1b9c; 12'hb08: x = 16'h1b98; 12'hb09: x = 16'h1b95; 12'hb0a: x = 16'h1b91; 12'hb0b: x = 16'h1b8e; 12'hb0c: x = 16'h1b8b; 12'hb0d: x = 16'h1b87; 12'hb0e: x = 16'h1b84; 12'hb0f: x = 16'h1b81; 12'hb10: x = 16'h1b7d; 12'hb11: x = 16'h1b7a; 12'hb12: x = 16'h1b77; 12'hb13: x = 16'h1b73; 12'hb14: x = 16'h1b70; 12'hb15: x = 16'h1b6c; 12'hb16: x = 16'h1b69; 12'hb17: x = 16'h1b66; 12'hb18: x = 16'h1b62; 12'hb19: x = 16'h1b5f; 12'hb1a: x = 16'h1b5c; 12'hb1b: x = 16'h1b58; 12'hb1c: x = 16'h1b55; 12'hb1d: x = 16'h1b51; 12'hb1e: x = 16'h1b4e; 12'hb1f: x = 16'h1b4b; 12'hb20: x = 16'h1b47; 12'hb21: x = 16'h1b44; 12'hb22: x = 16'h1b41; 12'hb23: x = 16'h1b3d; 12'hb24: x = 16'h1b3a; 12'hb25: x = 16'h1b36; 12'hb26: x = 16'h1b33; 12'hb27: x = 16'h1b30; 12'hb28: x = 16'h1b2c; 12'hb29: x = 16'h1b29; 12'hb2a: x = 16'h1b26; 12'hb2b: x = 16'h1b22; 12'hb2c: x = 16'h1b1f; 12'hb2d: x = 16'h1b1b; 12'hb2e: x = 16'h1b18; 12'hb2f: x = 16'h1b15; 12'hb30: x = 16'h1b11; 12'hb31: x = 16'h1b0e; 12'hb32: x = 16'h1b0b; 12'hb33: x = 16'h1b07; 12'hb34: x = 16'h1b04; 12'hb35: x = 16'h1b00; 12'hb36: x = 16'h1afd; 12'hb37: x = 16'h1afa; 12'hb38: x = 16'h1af6; 12'hb39: x = 16'h1af3; 12'hb3a: x = 16'h1aef; 12'hb3b: x = 16'h1aec; 12'hb3c: x = 16'h1ae9; 12'hb3d: x = 16'h1ae5; 12'hb3e: x = 16'h1ae2; 12'hb3f: x = 16'h1adf; 12'hb40: x = 16'h1adb; 12'hb41: x = 16'h1ad8; 12'hb42: x = 16'h1ad4; 12'hb43: x = 16'h1ad1; 12'hb44: x = 16'h1ace; 12'hb45: x = 16'h1aca; 12'hb46: x = 16'h1ac7; 12'hb47: x = 16'h1ac3; 12'hb48: x = 16'h1ac0; 12'hb49: x = 16'h1abd; 12'hb4a: x = 16'h1ab9; 12'hb4b: x = 16'h1ab6; 12'hb4c: x = 16'h1ab2; 12'hb4d: x = 16'h1aaf; 12'hb4e: x = 16'h1aac; 12'hb4f: x = 16'h1aa8; 12'hb50: x = 16'h1aa5; 12'hb51: x = 16'h1aa1; 12'hb52: x = 16'h1a9e; 12'hb53: x = 16'h1a9b; 12'hb54: x = 16'h1a97; 12'hb55: x = 16'h1a94; 12'hb56: x = 16'h1a90; 12'hb57: x = 16'h1a8d; 12'hb58: x = 16'h1a8a; 12'hb59: x = 16'h1a86; 12'hb5a: x = 16'h1a83; 12'hb5b: x = 16'h1a7f; 12'hb5c: x = 16'h1a7c; 12'hb5d: x = 16'h1a79; 12'hb5e: x = 16'h1a75; 12'hb5f: x = 16'h1a72; 12'hb60: x = 16'h1a6e; 12'hb61: x = 16'h1a6b; 12'hb62: x = 16'h1a68; 12'hb63: x = 16'h1a64; 12'hb64: x = 16'h1a61; 12'hb65: x = 16'h1a5d; 12'hb66: x = 16'h1a5a; 12'hb67: x = 16'h1a57; 12'hb68: x = 16'h1a53; 12'hb69: x = 16'h1a50; 12'hb6a: x = 16'h1a4c; 12'hb6b: x = 16'h1a49; 12'hb6c: x = 16'h1a46; 12'hb6d: x = 16'h1a42; 12'hb6e: x = 16'h1a3f; 12'hb6f: x = 16'h1a3b; 12'hb70: x = 16'h1a38; 12'hb71: x = 16'h1a34; 12'hb72: x = 16'h1a31; 12'hb73: x = 16'h1a2e; 12'hb74: x = 16'h1a2a; 12'hb75: x = 16'h1a27; 12'hb76: x = 16'h1a23; 12'hb77: x = 16'h1a20; 12'hb78: x = 16'h1a1d; 12'hb79: x = 16'h1a19; 12'hb7a: x = 16'h1a16; 12'hb7b: x = 16'h1a12; 12'hb7c: x = 16'h1a0f; 12'hb7d: x = 16'h1a0b; 12'hb7e: x = 16'h1a08; 12'hb7f: x = 16'h1a05; 12'hb80: x = 16'h1a01; 12'hb81: x = 16'h19fe; 12'hb82: x = 16'h19fa; 12'hb83: x = 16'h19f7; 12'hb84: x = 16'h19f3; 12'hb85: x = 16'h19f0; 12'hb86: x = 16'h19ed; 12'hb87: x = 16'h19e9; 12'hb88: x = 16'h19e6; 12'hb89: x = 16'h19e2; 12'hb8a: x = 16'h19df; 12'hb8b: x = 16'h19db; 12'hb8c: x = 16'h19d8; 12'hb8d: x = 16'h19d5; 12'hb8e: x = 16'h19d1; 12'hb8f: x = 16'h19ce; 12'hb90: x = 16'h19ca; 12'hb91: x = 16'h19c7; 12'hb92: x = 16'h19c3; 12'hb93: x = 16'h19c0; 12'hb94: x = 16'h19bd; 12'hb95: x = 16'h19b9; 12'hb96: x = 16'h19b6; 12'hb97: x = 16'h19b2; 12'hb98: x = 16'h19af; 12'hb99: x = 16'h19ab; 12'hb9a: x = 16'h19a8; 12'hb9b: x = 16'h19a4; 12'hb9c: x = 16'h19a1; 12'hb9d: x = 16'h199e; 12'hb9e: x = 16'h199a; 12'hb9f: x = 16'h1997; 12'hba0: x = 16'h1993; 12'hba1: x = 16'h1990; 12'hba2: x = 16'h198c; 12'hba3: x = 16'h1989; 12'hba4: x = 16'h1985; 12'hba5: x = 16'h1982; 12'hba6: x = 16'h197f; 12'hba7: x = 16'h197b; 12'hba8: x = 16'h1978; 12'hba9: x = 16'h1974; 12'hbaa: x = 16'h1971; 12'hbab: x = 16'h196d; 12'hbac: x = 16'h196a; 12'hbad: x = 16'h1966; 12'hbae: x = 16'h1963; 12'hbaf: x = 16'h1960; 12'hbb0: x = 16'h195c; 12'hbb1: x = 16'h1959; 12'hbb2: x = 16'h1955; 12'hbb3: x = 16'h1952; 12'hbb4: x = 16'h194e; 12'hbb5: x = 16'h194b; 12'hbb6: x = 16'h1947; 12'hbb7: x = 16'h1944; 12'hbb8: x = 16'h1940; 12'hbb9: x = 16'h193d; 12'hbba: x = 16'h1939; 12'hbbb: x = 16'h1936; 12'hbbc: x = 16'h1933; 12'hbbd: x = 16'h192f; 12'hbbe: x = 16'h192c; 12'hbbf: x = 16'h1928; 12'hbc0: x = 16'h1925; 12'hbc1: x = 16'h1921; 12'hbc2: x = 16'h191e; 12'hbc3: x = 16'h191a; 12'hbc4: x = 16'h1917; 12'hbc5: x = 16'h1913; 12'hbc6: x = 16'h1910; 12'hbc7: x = 16'h190c; 12'hbc8: x = 16'h1909; 12'hbc9: x = 16'h1905; 12'hbca: x = 16'h1902; 12'hbcb: x = 16'h18ff; 12'hbcc: x = 16'h18fb; 12'hbcd: x = 16'h18f8; 12'hbce: x = 16'h18f4; 12'hbcf: x = 16'h18f1; 12'hbd0: x = 16'h18ed; 12'hbd1: x = 16'h18ea; 12'hbd2: x = 16'h18e6; 12'hbd3: x = 16'h18e3; 12'hbd4: x = 16'h18df; 12'hbd5: x = 16'h18dc; 12'hbd6: x = 16'h18d8; 12'hbd7: x = 16'h18d5; 12'hbd8: x = 16'h18d1; 12'hbd9: x = 16'h18ce; 12'hbda: x = 16'h18ca; 12'hbdb: x = 16'h18c7; 12'hbdc: x = 16'h18c3; 12'hbdd: x = 16'h18c0; 12'hbde: x = 16'h18bc; 12'hbdf: x = 16'h18b9; 12'hbe0: x = 16'h18b5; 12'hbe1: x = 16'h18b2; 12'hbe2: x = 16'h18ae; 12'hbe3: x = 16'h18ab; 12'hbe4: x = 16'h18a7; 12'hbe5: x = 16'h18a4; 12'hbe6: x = 16'h18a0; 12'hbe7: x = 16'h189d; 12'hbe8: x = 16'h1899; 12'hbe9: x = 16'h1896; 12'hbea: x = 16'h1893; 12'hbeb: x = 16'h188f; 12'hbec: x = 16'h188c; 12'hbed: x = 16'h1888; 12'hbee: x = 16'h1885; 12'hbef: x = 16'h1881; 12'hbf0: x = 16'h187e; 12'hbf1: x = 16'h187a; 12'hbf2: x = 16'h1876; 12'hbf3: x = 16'h1873; 12'hbf4: x = 16'h186f; 12'hbf5: x = 16'h186c; 12'hbf6: x = 16'h1868; 12'hbf7: x = 16'h1865; 12'hbf8: x = 16'h1861; 12'hbf9: x = 16'h185e; 12'hbfa: x = 16'h185a; 12'hbfb: x = 16'h1857; 12'hbfc: x = 16'h1853; 12'hbfd: x = 16'h1850; 12'hbfe: x = 16'h184c; 12'hbff: x = 16'h1849; 12'hc00: x = 16'h1845; 12'hc01: x = 16'h1842; 12'hc02: x = 16'h183e; 12'hc03: x = 16'h183b; 12'hc04: x = 16'h1837; 12'hc05: x = 16'h1834; 12'hc06: x = 16'h1830; 12'hc07: x = 16'h182d; 12'hc08: x = 16'h1829; 12'hc09: x = 16'h1826; 12'hc0a: x = 16'h1822; 12'hc0b: x = 16'h181f; 12'hc0c: x = 16'h181b; 12'hc0d: x = 16'h1818; 12'hc0e: x = 16'h1814; 12'hc0f: x = 16'h1811; 12'hc10: x = 16'h180d; 12'hc11: x = 16'h1809; 12'hc12: x = 16'h1806; 12'hc13: x = 16'h1802; 12'hc14: x = 16'h17ff; 12'hc15: x = 16'h17fb; 12'hc16: x = 16'h17f8; 12'hc17: x = 16'h17f4; 12'hc18: x = 16'h17f1; 12'hc19: x = 16'h17ed; 12'hc1a: x = 16'h17ea; 12'hc1b: x = 16'h17e6; 12'hc1c: x = 16'h17e3; 12'hc1d: x = 16'h17df; 12'hc1e: x = 16'h17dc; 12'hc1f: x = 16'h17d8; 12'hc20: x = 16'h17d4; 12'hc21: x = 16'h17d1; 12'hc22: x = 16'h17cd; 12'hc23: x = 16'h17ca; 12'hc24: x = 16'h17c6; 12'hc25: x = 16'h17c3; 12'hc26: x = 16'h17bf; 12'hc27: x = 16'h17bc; 12'hc28: x = 16'h17b8; 12'hc29: x = 16'h17b4; 12'hc2a: x = 16'h17b1; 12'hc2b: x = 16'h17ad; 12'hc2c: x = 16'h17aa; 12'hc2d: x = 16'h17a6; 12'hc2e: x = 16'h17a3; 12'hc2f: x = 16'h179f; 12'hc30: x = 16'h179c; 12'hc31: x = 16'h1798; 12'hc32: x = 16'h1794; 12'hc33: x = 16'h1791; 12'hc34: x = 16'h178d; 12'hc35: x = 16'h178a; 12'hc36: x = 16'h1786; 12'hc37: x = 16'h1783; 12'hc38: x = 16'h177f; 12'hc39: x = 16'h177c; 12'hc3a: x = 16'h1778; 12'hc3b: x = 16'h1774; 12'hc3c: x = 16'h1771; 12'hc3d: x = 16'h176d; 12'hc3e: x = 16'h176a; 12'hc3f: x = 16'h1766; 12'hc40: x = 16'h1763; 12'hc41: x = 16'h175f; 12'hc42: x = 16'h175b; 12'hc43: x = 16'h1758; 12'hc44: x = 16'h1754; 12'hc45: x = 16'h1751; 12'hc46: x = 16'h174d; 12'hc47: x = 16'h1749; 12'hc48: x = 16'h1746; 12'hc49: x = 16'h1742; 12'hc4a: x = 16'h173f; 12'hc4b: x = 16'h173b; 12'hc4c: x = 16'h1738; 12'hc4d: x = 16'h1734; 12'hc4e: x = 16'h1730; 12'hc4f: x = 16'h172d; 12'hc50: x = 16'h1729; 12'hc51: x = 16'h1726; 12'hc52: x = 16'h1722; 12'hc53: x = 16'h171e; 12'hc54: x = 16'h171b; 12'hc55: x = 16'h1717; 12'hc56: x = 16'h1714; 12'hc57: x = 16'h1710; 12'hc58: x = 16'h170c; 12'hc59: x = 16'h1709; 12'hc5a: x = 16'h1705; 12'hc5b: x = 16'h1702; 12'hc5c: x = 16'h16fe; 12'hc5d: x = 16'h16fa; 12'hc5e: x = 16'h16f7; 12'hc5f: x = 16'h16f3; 12'hc60: x = 16'h16f0; 12'hc61: x = 16'h16ec; 12'hc62: x = 16'h16e8; 12'hc63: x = 16'h16e5; 12'hc64: x = 16'h16e1; 12'hc65: x = 16'h16de; 12'hc66: x = 16'h16da; 12'hc67: x = 16'h16d6; 12'hc68: x = 16'h16d3; 12'hc69: x = 16'h16cf; 12'hc6a: x = 16'h16cc; 12'hc6b: x = 16'h16c8; 12'hc6c: x = 16'h16c4; 12'hc6d: x = 16'h16c1; 12'hc6e: x = 16'h16bd; 12'hc6f: x = 16'h16b9; 12'hc70: x = 16'h16b6; 12'hc71: x = 16'h16b2; 12'hc72: x = 16'h16af; 12'hc73: x = 16'h16ab; 12'hc74: x = 16'h16a7; 12'hc75: x = 16'h16a4; 12'hc76: x = 16'h16a0; 12'hc77: x = 16'h169c; 12'hc78: x = 16'h1699; 12'hc79: x = 16'h1695; 12'hc7a: x = 16'h1691; 12'hc7b: x = 16'h168e; 12'hc7c: x = 16'h168a; 12'hc7d: x = 16'h1687; 12'hc7e: x = 16'h1683; 12'hc7f: x = 16'h167f; 12'hc80: x = 16'h167c; 12'hc81: x = 16'h1678; 12'hc82: x = 16'h1674; 12'hc83: x = 16'h1671; 12'hc84: x = 16'h166d; 12'hc85: x = 16'h1669; 12'hc86: x = 16'h1666; 12'hc87: x = 16'h1662; 12'hc88: x = 16'h165e; 12'hc89: x = 16'h165b; 12'hc8a: x = 16'h1657; 12'hc8b: x = 16'h1653; 12'hc8c: x = 16'h1650; 12'hc8d: x = 16'h164c; 12'hc8e: x = 16'h1649; 12'hc8f: x = 16'h1645; 12'hc90: x = 16'h1641; 12'hc91: x = 16'h163e; 12'hc92: x = 16'h163a; 12'hc93: x = 16'h1636; 12'hc94: x = 16'h1633; 12'hc95: x = 16'h162f; 12'hc96: x = 16'h162b; 12'hc97: x = 16'h1628; 12'hc98: x = 16'h1624; 12'hc99: x = 16'h1620; 12'hc9a: x = 16'h161c; 12'hc9b: x = 16'h1619; 12'hc9c: x = 16'h1615; 12'hc9d: x = 16'h1611; 12'hc9e: x = 16'h160e; 12'hc9f: x = 16'h160a; 12'hca0: x = 16'h1606; 12'hca1: x = 16'h1603; 12'hca2: x = 16'h15ff; 12'hca3: x = 16'h15fb; 12'hca4: x = 16'h15f8; 12'hca5: x = 16'h15f4; 12'hca6: x = 16'h15f0; 12'hca7: x = 16'h15ed; 12'hca8: x = 16'h15e9; 12'hca9: x = 16'h15e5; 12'hcaa: x = 16'h15e2; 12'hcab: x = 16'h15de; 12'hcac: x = 16'h15da; 12'hcad: x = 16'h15d6; 12'hcae: x = 16'h15d3; 12'hcaf: x = 16'h15cf; 12'hcb0: x = 16'h15cb; 12'hcb1: x = 16'h15c8; 12'hcb2: x = 16'h15c4; 12'hcb3: x = 16'h15c0; 12'hcb4: x = 16'h15bd; 12'hcb5: x = 16'h15b9; 12'hcb6: x = 16'h15b5; 12'hcb7: x = 16'h15b1; 12'hcb8: x = 16'h15ae; 12'hcb9: x = 16'h15aa; 12'hcba: x = 16'h15a6; 12'hcbb: x = 16'h15a3; 12'hcbc: x = 16'h159f; 12'hcbd: x = 16'h159b; 12'hcbe: x = 16'h1597; 12'hcbf: x = 16'h1594; 12'hcc0: x = 16'h1590; 12'hcc1: x = 16'h158c; 12'hcc2: x = 16'h1588; 12'hcc3: x = 16'h1585; 12'hcc4: x = 16'h1581; 12'hcc5: x = 16'h157d; 12'hcc6: x = 16'h157a; 12'hcc7: x = 16'h1576; 12'hcc8: x = 16'h1572; 12'hcc9: x = 16'h156e; 12'hcca: x = 16'h156b; 12'hccb: x = 16'h1567; 12'hccc: x = 16'h1563; 12'hccd: x = 16'h155f; 12'hcce: x = 16'h155c; 12'hccf: x = 16'h1558; 12'hcd0: x = 16'h1554; 12'hcd1: x = 16'h1550; 12'hcd2: x = 16'h154d; 12'hcd3: x = 16'h1549; 12'hcd4: x = 16'h1545; 12'hcd5: x = 16'h1541; 12'hcd6: x = 16'h153e; 12'hcd7: x = 16'h153a; 12'hcd8: x = 16'h1536; 12'hcd9: x = 16'h1532; 12'hcda: x = 16'h152f; 12'hcdb: x = 16'h152b; 12'hcdc: x = 16'h1527; 12'hcdd: x = 16'h1523; 12'hcde: x = 16'h1520; 12'hcdf: x = 16'h151c; 12'hce0: x = 16'h1518; 12'hce1: x = 16'h1514; 12'hce2: x = 16'h1510; 12'hce3: x = 16'h150d; 12'hce4: x = 16'h1509; 12'hce5: x = 16'h1505; 12'hce6: x = 16'h1501; 12'hce7: x = 16'h14fe; 12'hce8: x = 16'h14fa; 12'hce9: x = 16'h14f6; 12'hcea: x = 16'h14f2; 12'hceb: x = 16'h14ee; 12'hcec: x = 16'h14eb; 12'hced: x = 16'h14e7; 12'hcee: x = 16'h14e3; 12'hcef: x = 16'h14df; 12'hcf0: x = 16'h14dc; 12'hcf1: x = 16'h14d8; 12'hcf2: x = 16'h14d4; 12'hcf3: x = 16'h14d0; 12'hcf4: x = 16'h14cc; 12'hcf5: x = 16'h14c9; 12'hcf6: x = 16'h14c5; 12'hcf7: x = 16'h14c1; 12'hcf8: x = 16'h14bd; 12'hcf9: x = 16'h14b9; 12'hcfa: x = 16'h14b5; 12'hcfb: x = 16'h14b2; 12'hcfc: x = 16'h14ae; 12'hcfd: x = 16'h14aa; 12'hcfe: x = 16'h14a6; 12'hcff: x = 16'h14a2; 12'hd00: x = 16'h149f; 12'hd01: x = 16'h149b; 12'hd02: x = 16'h1497; 12'hd03: x = 16'h1493; 12'hd04: x = 16'h148f; 12'hd05: x = 16'h148b; 12'hd06: x = 16'h1488; 12'hd07: x = 16'h1484; 12'hd08: x = 16'h1480; 12'hd09: x = 16'h147c; 12'hd0a: x = 16'h1478; 12'hd0b: x = 16'h1474; 12'hd0c: x = 16'h1471; 12'hd0d: x = 16'h146d; 12'hd0e: x = 16'h1469; 12'hd0f: x = 16'h1465; 12'hd10: x = 16'h1461; 12'hd11: x = 16'h145d; 12'hd12: x = 16'h145a; 12'hd13: x = 16'h1456; 12'hd14: x = 16'h1452; 12'hd15: x = 16'h144e; 12'hd16: x = 16'h144a; 12'hd17: x = 16'h1446; 12'hd18: x = 16'h1442; 12'hd19: x = 16'h143f; 12'hd1a: x = 16'h143b; 12'hd1b: x = 16'h1437; 12'hd1c: x = 16'h1433; 12'hd1d: x = 16'h142f; 12'hd1e: x = 16'h142b; 12'hd1f: x = 16'h1427; 12'hd20: x = 16'h1424; 12'hd21: x = 16'h1420; 12'hd22: x = 16'h141c; 12'hd23: x = 16'h1418; 12'hd24: x = 16'h1414; 12'hd25: x = 16'h1410; 12'hd26: x = 16'h140c; 12'hd27: x = 16'h1408; 12'hd28: x = 16'h1404; 12'hd29: x = 16'h1401; 12'hd2a: x = 16'h13fd; 12'hd2b: x = 16'h13f9; 12'hd2c: x = 16'h13f5; 12'hd2d: x = 16'h13f1; 12'hd2e: x = 16'h13ed; 12'hd2f: x = 16'h13e9; 12'hd30: x = 16'h13e5; 12'hd31: x = 16'h13e1; 12'hd32: x = 16'h13dd; 12'hd33: x = 16'h13da; 12'hd34: x = 16'h13d6; 12'hd35: x = 16'h13d2; 12'hd36: x = 16'h13ce; 12'hd37: x = 16'h13ca; 12'hd38: x = 16'h13c6; 12'hd39: x = 16'h13c2; 12'hd3a: x = 16'h13be; 12'hd3b: x = 16'h13ba; 12'hd3c: x = 16'h13b6; 12'hd3d: x = 16'h13b2; 12'hd3e: x = 16'h13ae; 12'hd3f: x = 16'h13ab; 12'hd40: x = 16'h13a7; 12'hd41: x = 16'h13a3; 12'hd42: x = 16'h139f; 12'hd43: x = 16'h139b; 12'hd44: x = 16'h1397; 12'hd45: x = 16'h1393; 12'hd46: x = 16'h138f; 12'hd47: x = 16'h138b; 12'hd48: x = 16'h1387; 12'hd49: x = 16'h1383; 12'hd4a: x = 16'h137f; 12'hd4b: x = 16'h137b; 12'hd4c: x = 16'h1377; 12'hd4d: x = 16'h1373; 12'hd4e: x = 16'h136f; 12'hd4f: x = 16'h136b; 12'hd50: x = 16'h1367; 12'hd51: x = 16'h1363; 12'hd52: x = 16'h1360; 12'hd53: x = 16'h135c; 12'hd54: x = 16'h1358; 12'hd55: x = 16'h1354; 12'hd56: x = 16'h1350; 12'hd57: x = 16'h134c; 12'hd58: x = 16'h1348; 12'hd59: x = 16'h1344; 12'hd5a: x = 16'h1340; 12'hd5b: x = 16'h133c; 12'hd5c: x = 16'h1338; 12'hd5d: x = 16'h1334; 12'hd5e: x = 16'h1330; 12'hd5f: x = 16'h132c; 12'hd60: x = 16'h1328; 12'hd61: x = 16'h1324; 12'hd62: x = 16'h1320; 12'hd63: x = 16'h131c; 12'hd64: x = 16'h1318; 12'hd65: x = 16'h1314; 12'hd66: x = 16'h1310; 12'hd67: x = 16'h130c; 12'hd68: x = 16'h1308; 12'hd69: x = 16'h1304; 12'hd6a: x = 16'h1300; 12'hd6b: x = 16'h12fc; 12'hd6c: x = 16'h12f8; 12'hd6d: x = 16'h12f4; 12'hd6e: x = 16'h12f0; 12'hd6f: x = 16'h12ec; 12'hd70: x = 16'h12e8; 12'hd71: x = 16'h12e4; 12'hd72: x = 16'h12e0; 12'hd73: x = 16'h12db; 12'hd74: x = 16'h12d7; 12'hd75: x = 16'h12d3; 12'hd76: x = 16'h12cf; 12'hd77: x = 16'h12cb; 12'hd78: x = 16'h12c7; 12'hd79: x = 16'h12c3; 12'hd7a: x = 16'h12bf; 12'hd7b: x = 16'h12bb; 12'hd7c: x = 16'h12b7; 12'hd7d: x = 16'h12b3; 12'hd7e: x = 16'h12af; 12'hd7f: x = 16'h12ab; 12'hd80: x = 16'h12a7; 12'hd81: x = 16'h12a3; 12'hd82: x = 16'h129f; 12'hd83: x = 16'h129b; 12'hd84: x = 16'h1297; 12'hd85: x = 16'h1292; 12'hd86: x = 16'h128e; 12'hd87: x = 16'h128a; 12'hd88: x = 16'h1286; 12'hd89: x = 16'h1282; 12'hd8a: x = 16'h127e; 12'hd8b: x = 16'h127a; 12'hd8c: x = 16'h1276; 12'hd8d: x = 16'h1272; 12'hd8e: x = 16'h126e; 12'hd8f: x = 16'h126a; 12'hd90: x = 16'h1265; 12'hd91: x = 16'h1261; 12'hd92: x = 16'h125d; 12'hd93: x = 16'h1259; 12'hd94: x = 16'h1255; 12'hd95: x = 16'h1251; 12'hd96: x = 16'h124d; 12'hd97: x = 16'h1249; 12'hd98: x = 16'h1245; 12'hd99: x = 16'h1240; 12'hd9a: x = 16'h123c; 12'hd9b: x = 16'h1238; 12'hd9c: x = 16'h1234; 12'hd9d: x = 16'h1230; 12'hd9e: x = 16'h122c; 12'hd9f: x = 16'h1228; 12'hda0: x = 16'h1223; 12'hda1: x = 16'h121f; 12'hda2: x = 16'h121b; 12'hda3: x = 16'h1217; 12'hda4: x = 16'h1213; 12'hda5: x = 16'h120f; 12'hda6: x = 16'h120b; 12'hda7: x = 16'h1206; 12'hda8: x = 16'h1202; 12'hda9: x = 16'h11fe; 12'hdaa: x = 16'h11fa; 12'hdab: x = 16'h11f6; 12'hdac: x = 16'h11f2; 12'hdad: x = 16'h11ed; 12'hdae: x = 16'h11e9; 12'hdaf: x = 16'h11e5; 12'hdb0: x = 16'h11e1; 12'hdb1: x = 16'h11dd; 12'hdb2: x = 16'h11d8; 12'hdb3: x = 16'h11d4; 12'hdb4: x = 16'h11d0; 12'hdb5: x = 16'h11cc; 12'hdb6: x = 16'h11c8; 12'hdb7: x = 16'h11c3; 12'hdb8: x = 16'h11bf; 12'hdb9: x = 16'h11bb; 12'hdba: x = 16'h11b7; 12'hdbb: x = 16'h11b3; 12'hdbc: x = 16'h11ae; 12'hdbd: x = 16'h11aa; 12'hdbe: x = 16'h11a6; 12'hdbf: x = 16'h11a2; 12'hdc0: x = 16'h119e; 12'hdc1: x = 16'h1199; 12'hdc2: x = 16'h1195; 12'hdc3: x = 16'h1191; 12'hdc4: x = 16'h118d; 12'hdc5: x = 16'h1188; 12'hdc6: x = 16'h1184; 12'hdc7: x = 16'h1180; 12'hdc8: x = 16'h117c; 12'hdc9: x = 16'h1177; 12'hdca: x = 16'h1173; 12'hdcb: x = 16'h116f; 12'hdcc: x = 16'h116b; 12'hdcd: x = 16'h1166; 12'hdce: x = 16'h1162; 12'hdcf: x = 16'h115e; 12'hdd0: x = 16'h115a; 12'hdd1: x = 16'h1155; 12'hdd2: x = 16'h1151; 12'hdd3: x = 16'h114d; 12'hdd4: x = 16'h1148; 12'hdd5: x = 16'h1144; 12'hdd6: x = 16'h1140; 12'hdd7: x = 16'h113c; 12'hdd8: x = 16'h1137; 12'hdd9: x = 16'h1133; 12'hdda: x = 16'h112f; 12'hddb: x = 16'h112a; 12'hddc: x = 16'h1126; 12'hddd: x = 16'h1122; 12'hdde: x = 16'h111d; 12'hddf: x = 16'h1119; 12'hde0: x = 16'h1115; 12'hde1: x = 16'h1111; 12'hde2: x = 16'h110c; 12'hde3: x = 16'h1108; 12'hde4: x = 16'h1104; 12'hde5: x = 16'h10ff; 12'hde6: x = 16'h10fb; 12'hde7: x = 16'h10f7; 12'hde8: x = 16'h10f2; 12'hde9: x = 16'h10ee; 12'hdea: x = 16'h10e9; 12'hdeb: x = 16'h10e5; 12'hdec: x = 16'h10e1; 12'hded: x = 16'h10dc; 12'hdee: x = 16'h10d8; 12'hdef: x = 16'h10d4; 12'hdf0: x = 16'h10cf; 12'hdf1: x = 16'h10cb; 12'hdf2: x = 16'h10c7; 12'hdf3: x = 16'h10c2; 12'hdf4: x = 16'h10be; 12'hdf5: x = 16'h10b9; 12'hdf6: x = 16'h10b5; 12'hdf7: x = 16'h10b1; 12'hdf8: x = 16'h10ac; 12'hdf9: x = 16'h10a8; 12'hdfa: x = 16'h10a3; 12'hdfb: x = 16'h109f; 12'hdfc: x = 16'h109b; 12'hdfd: x = 16'h1096; 12'hdfe: x = 16'h1092; 12'hdff: x = 16'h108d; 12'he00: x = 16'h1089; 12'he01: x = 16'h1085; 12'he02: x = 16'h1080; 12'he03: x = 16'h107c; 12'he04: x = 16'h1077; 12'he05: x = 16'h1073; 12'he06: x = 16'h106e; 12'he07: x = 16'h106a; 12'he08: x = 16'h1065; 12'he09: x = 16'h1061; 12'he0a: x = 16'h105d; 12'he0b: x = 16'h1058; 12'he0c: x = 16'h1054; 12'he0d: x = 16'h104f; 12'he0e: x = 16'h104b; 12'he0f: x = 16'h1046; 12'he10: x = 16'h1042; 12'he11: x = 16'h103d; 12'he12: x = 16'h1039; 12'he13: x = 16'h1034; 12'he14: x = 16'h1030; 12'he15: x = 16'h102b; 12'he16: x = 16'h1027; 12'he17: x = 16'h1022; 12'he18: x = 16'h101e; 12'he19: x = 16'h1019; 12'he1a: x = 16'h1015; 12'he1b: x = 16'h1010; 12'he1c: x = 16'h100c; 12'he1d: x = 16'h1007; 12'he1e: x = 16'h1003; 12'he1f: x = 16'h ffe; 12'he20: x = 16'h ffa; 12'he21: x = 16'h ff5; 12'he22: x = 16'h ff1; 12'he23: x = 16'h fec; 12'he24: x = 16'h fe7; 12'he25: x = 16'h fe3; 12'he26: x = 16'h fde; 12'he27: x = 16'h fda; 12'he28: x = 16'h fd5; 12'he29: x = 16'h fd1; 12'he2a: x = 16'h fcc; 12'he2b: x = 16'h fc7; 12'he2c: x = 16'h fc3; 12'he2d: x = 16'h fbe; 12'he2e: x = 16'h fba; 12'he2f: x = 16'h fb5; 12'he30: x = 16'h fb1; 12'he31: x = 16'h fac; 12'he32: x = 16'h fa7; 12'he33: x = 16'h fa3; 12'he34: x = 16'h f9e; 12'he35: x = 16'h f99; 12'he36: x = 16'h f95; 12'he37: x = 16'h f90; 12'he38: x = 16'h f8c; 12'he39: x = 16'h f87; 12'he3a: x = 16'h f82; 12'he3b: x = 16'h f7e; 12'he3c: x = 16'h f79; 12'he3d: x = 16'h f74; 12'he3e: x = 16'h f70; 12'he3f: x = 16'h f6b; 12'he40: x = 16'h f66; 12'he41: x = 16'h f62; 12'he42: x = 16'h f5d; 12'he43: x = 16'h f58; 12'he44: x = 16'h f54; 12'he45: x = 16'h f4f; 12'he46: x = 16'h f4a; 12'he47: x = 16'h f46; 12'he48: x = 16'h f41; 12'he49: x = 16'h f3c; 12'he4a: x = 16'h f38; 12'he4b: x = 16'h f33; 12'he4c: x = 16'h f2e; 12'he4d: x = 16'h f29; 12'he4e: x = 16'h f25; 12'he4f: x = 16'h f20; 12'he50: x = 16'h f1b; 12'he51: x = 16'h f16; 12'he52: x = 16'h f12; 12'he53: x = 16'h f0d; 12'he54: x = 16'h f08; 12'he55: x = 16'h f03; 12'he56: x = 16'h eff; 12'he57: x = 16'h efa; 12'he58: x = 16'h ef5; 12'he59: x = 16'h ef0; 12'he5a: x = 16'h eec; 12'he5b: x = 16'h ee7; 12'he5c: x = 16'h ee2; 12'he5d: x = 16'h edd; 12'he5e: x = 16'h ed8; 12'he5f: x = 16'h ed4; 12'he60: x = 16'h ecf; 12'he61: x = 16'h eca; 12'he62: x = 16'h ec5; 12'he63: x = 16'h ec0; 12'he64: x = 16'h ebc; 12'he65: x = 16'h eb7; 12'he66: x = 16'h eb2; 12'he67: x = 16'h ead; 12'he68: x = 16'h ea8; 12'he69: x = 16'h ea3; 12'he6a: x = 16'h e9f; 12'he6b: x = 16'h e9a; 12'he6c: x = 16'h e95; 12'he6d: x = 16'h e90; 12'he6e: x = 16'h e8b; 12'he6f: x = 16'h e86; 12'he70: x = 16'h e81; 12'he71: x = 16'h e7c; 12'he72: x = 16'h e77; 12'he73: x = 16'h e73; 12'he74: x = 16'h e6e; 12'he75: x = 16'h e69; 12'he76: x = 16'h e64; 12'he77: x = 16'h e5f; 12'he78: x = 16'h e5a; 12'he79: x = 16'h e55; 12'he7a: x = 16'h e50; 12'he7b: x = 16'h e4b; 12'he7c: x = 16'h e46; 12'he7d: x = 16'h e41; 12'he7e: x = 16'h e3c; 12'he7f: x = 16'h e37; 12'he80: x = 16'h e32; 12'he81: x = 16'h e2d; 12'he82: x = 16'h e28; 12'he83: x = 16'h e23; 12'he84: x = 16'h e1e; 12'he85: x = 16'h e19; 12'he86: x = 16'h e14; 12'he87: x = 16'h e0f; 12'he88: x = 16'h e0a; 12'he89: x = 16'h e05; 12'he8a: x = 16'h e00; 12'he8b: x = 16'h dfb; 12'he8c: x = 16'h df6; 12'he8d: x = 16'h df1; 12'he8e: x = 16'h dec; 12'he8f: x = 16'h de7; 12'he90: x = 16'h de2; 12'he91: x = 16'h ddd; 12'he92: x = 16'h dd8; 12'he93: x = 16'h dd3; 12'he94: x = 16'h dce; 12'he95: x = 16'h dc9; 12'he96: x = 16'h dc4; 12'he97: x = 16'h dbe; 12'he98: x = 16'h db9; 12'he99: x = 16'h db4; 12'he9a: x = 16'h daf; 12'he9b: x = 16'h daa; 12'he9c: x = 16'h da5; 12'he9d: x = 16'h da0; 12'he9e: x = 16'h d9b; 12'he9f: x = 16'h d95; 12'hea0: x = 16'h d90; 12'hea1: x = 16'h d8b; 12'hea2: x = 16'h d86; 12'hea3: x = 16'h d81; 12'hea4: x = 16'h d7c; 12'hea5: x = 16'h d76; 12'hea6: x = 16'h d71; 12'hea7: x = 16'h d6c; 12'hea8: x = 16'h d67; 12'hea9: x = 16'h d62; 12'heaa: x = 16'h d5c; 12'heab: x = 16'h d57; 12'heac: x = 16'h d52; 12'head: x = 16'h d4d; 12'heae: x = 16'h d47; 12'heaf: x = 16'h d42; 12'heb0: x = 16'h d3d; 12'heb1: x = 16'h d38; 12'heb2: x = 16'h d32; 12'heb3: x = 16'h d2d; 12'heb4: x = 16'h d28; 12'heb5: x = 16'h d22; 12'heb6: x = 16'h d1d; 12'heb7: x = 16'h d18; 12'heb8: x = 16'h d13; 12'heb9: x = 16'h d0d; 12'heba: x = 16'h d08; 12'hebb: x = 16'h d03; 12'hebc: x = 16'h cfd; 12'hebd: x = 16'h cf8; 12'hebe: x = 16'h cf2; 12'hebf: x = 16'h ced; 12'hec0: x = 16'h ce8; 12'hec1: x = 16'h ce2; 12'hec2: x = 16'h cdd; 12'hec3: x = 16'h cd8; 12'hec4: x = 16'h cd2; 12'hec5: x = 16'h ccd; 12'hec6: x = 16'h cc7; 12'hec7: x = 16'h cc2; 12'hec8: x = 16'h cbc; 12'hec9: x = 16'h cb7; 12'heca: x = 16'h cb2; 12'hecb: x = 16'h cac; 12'hecc: x = 16'h ca7; 12'hecd: x = 16'h ca1; 12'hece: x = 16'h c9c; 12'hecf: x = 16'h c96; 12'hed0: x = 16'h c91; 12'hed1: x = 16'h c8b; 12'hed2: x = 16'h c86; 12'hed3: x = 16'h c80; 12'hed4: x = 16'h c7b; 12'hed5: x = 16'h c75; 12'hed6: x = 16'h c70; 12'hed7: x = 16'h c6a; 12'hed8: x = 16'h c64; 12'hed9: x = 16'h c5f; 12'heda: x = 16'h c59; 12'hedb: x = 16'h c54; 12'hedc: x = 16'h c4e; 12'hedd: x = 16'h c49; 12'hede: x = 16'h c43; 12'hedf: x = 16'h c3d; 12'hee0: x = 16'h c38; 12'hee1: x = 16'h c32; 12'hee2: x = 16'h c2c; 12'hee3: x = 16'h c27; 12'hee4: x = 16'h c21; 12'hee5: x = 16'h c1b; 12'hee6: x = 16'h c16; 12'hee7: x = 16'h c10; 12'hee8: x = 16'h c0a; 12'hee9: x = 16'h c05; 12'heea: x = 16'h bff; 12'heeb: x = 16'h bf9; 12'heec: x = 16'h bf3; 12'heed: x = 16'h bee; 12'heee: x = 16'h be8; 12'heef: x = 16'h be2; 12'hef0: x = 16'h bdc; 12'hef1: x = 16'h bd7; 12'hef2: x = 16'h bd1; 12'hef3: x = 16'h bcb; 12'hef4: x = 16'h bc5; 12'hef5: x = 16'h bbf; 12'hef6: x = 16'h bba; 12'hef7: x = 16'h bb4; 12'hef8: x = 16'h bae; 12'hef9: x = 16'h ba8; 12'hefa: x = 16'h ba2; 12'hefb: x = 16'h b9c; 12'hefc: x = 16'h b96; 12'hefd: x = 16'h b90; 12'hefe: x = 16'h b8b; 12'heff: x = 16'h b85; 12'hf00: x = 16'h b7f; 12'hf01: x = 16'h b79; 12'hf02: x = 16'h b73; 12'hf03: x = 16'h b6d; 12'hf04: x = 16'h b67; 12'hf05: x = 16'h b61; 12'hf06: x = 16'h b5b; 12'hf07: x = 16'h b55; 12'hf08: x = 16'h b4f; 12'hf09: x = 16'h b49; 12'hf0a: x = 16'h b43; 12'hf0b: x = 16'h b3d; 12'hf0c: x = 16'h b37; 12'hf0d: x = 16'h b31; 12'hf0e: x = 16'h b2a; 12'hf0f: x = 16'h b24; 12'hf10: x = 16'h b1e; 12'hf11: x = 16'h b18; 12'hf12: x = 16'h b12; 12'hf13: x = 16'h b0c; 12'hf14: x = 16'h b06; 12'hf15: x = 16'h b00; 12'hf16: x = 16'h af9; 12'hf17: x = 16'h af3; 12'hf18: x = 16'h aed; 12'hf19: x = 16'h ae7; 12'hf1a: x = 16'h ae1; 12'hf1b: x = 16'h ada; 12'hf1c: x = 16'h ad4; 12'hf1d: x = 16'h ace; 12'hf1e: x = 16'h ac8; 12'hf1f: x = 16'h ac1; 12'hf20: x = 16'h abb; 12'hf21: x = 16'h ab5; 12'hf22: x = 16'h aae; 12'hf23: x = 16'h aa8; 12'hf24: x = 16'h aa2; 12'hf25: x = 16'h a9b; 12'hf26: x = 16'h a95; 12'hf27: x = 16'h a8e; 12'hf28: x = 16'h a88; 12'hf29: x = 16'h a82; 12'hf2a: x = 16'h a7b; 12'hf2b: x = 16'h a75; 12'hf2c: x = 16'h a6e; 12'hf2d: x = 16'h a68; 12'hf2e: x = 16'h a61; 12'hf2f: x = 16'h a5b; 12'hf30: x = 16'h a54; 12'hf31: x = 16'h a4e; 12'hf32: x = 16'h a47; 12'hf33: x = 16'h a41; 12'hf34: x = 16'h a3a; 12'hf35: x = 16'h a33; 12'hf36: x = 16'h a2d; 12'hf37: x = 16'h a26; 12'hf38: x = 16'h a20; 12'hf39: x = 16'h a19; 12'hf3a: x = 16'h a12; 12'hf3b: x = 16'h a0c; 12'hf3c: x = 16'h a05; 12'hf3d: x = 16'h 9fe; 12'hf3e: x = 16'h 9f7; 12'hf3f: x = 16'h 9f1; 12'hf40: x = 16'h 9ea; 12'hf41: x = 16'h 9e3; 12'hf42: x = 16'h 9dc; 12'hf43: x = 16'h 9d6; 12'hf44: x = 16'h 9cf; 12'hf45: x = 16'h 9c8; 12'hf46: x = 16'h 9c1; 12'hf47: x = 16'h 9ba; 12'hf48: x = 16'h 9b3; 12'hf49: x = 16'h 9ac; 12'hf4a: x = 16'h 9a5; 12'hf4b: x = 16'h 99e; 12'hf4c: x = 16'h 997; 12'hf4d: x = 16'h 990; 12'hf4e: x = 16'h 989; 12'hf4f: x = 16'h 982; 12'hf50: x = 16'h 97b; 12'hf51: x = 16'h 974; 12'hf52: x = 16'h 96d; 12'hf53: x = 16'h 966; 12'hf54: x = 16'h 95f; 12'hf55: x = 16'h 958; 12'hf56: x = 16'h 951; 12'hf57: x = 16'h 94a; 12'hf58: x = 16'h 942; 12'hf59: x = 16'h 93b; 12'hf5a: x = 16'h 934; 12'hf5b: x = 16'h 92d; 12'hf5c: x = 16'h 925; 12'hf5d: x = 16'h 91e; 12'hf5e: x = 16'h 917; 12'hf5f: x = 16'h 90f; 12'hf60: x = 16'h 908; 12'hf61: x = 16'h 901; 12'hf62: x = 16'h 8f9; 12'hf63: x = 16'h 8f2; 12'hf64: x = 16'h 8ea; 12'hf65: x = 16'h 8e3; 12'hf66: x = 16'h 8db; 12'hf67: x = 16'h 8d4; 12'hf68: x = 16'h 8cc; 12'hf69: x = 16'h 8c5; 12'hf6a: x = 16'h 8bd; 12'hf6b: x = 16'h 8b6; 12'hf6c: x = 16'h 8ae; 12'hf6d: x = 16'h 8a6; 12'hf6e: x = 16'h 89f; 12'hf6f: x = 16'h 897; 12'hf70: x = 16'h 88f; 12'hf71: x = 16'h 887; 12'hf72: x = 16'h 880; 12'hf73: x = 16'h 878; 12'hf74: x = 16'h 870; 12'hf75: x = 16'h 868; 12'hf76: x = 16'h 860; 12'hf77: x = 16'h 858; 12'hf78: x = 16'h 850; 12'hf79: x = 16'h 848; 12'hf7a: x = 16'h 840; 12'hf7b: x = 16'h 838; 12'hf7c: x = 16'h 830; 12'hf7d: x = 16'h 828; 12'hf7e: x = 16'h 820; 12'hf7f: x = 16'h 818; 12'hf80: x = 16'h 810; 12'hf81: x = 16'h 808; 12'hf82: x = 16'h 7ff; 12'hf83: x = 16'h 7f7; 12'hf84: x = 16'h 7ef; 12'hf85: x = 16'h 7e6; 12'hf86: x = 16'h 7de; 12'hf87: x = 16'h 7d6; 12'hf88: x = 16'h 7cd; 12'hf89: x = 16'h 7c5; 12'hf8a: x = 16'h 7bc; 12'hf8b: x = 16'h 7b4; 12'hf8c: x = 16'h 7ab; 12'hf8d: x = 16'h 7a3; 12'hf8e: x = 16'h 79a; 12'hf8f: x = 16'h 791; 12'hf90: x = 16'h 789; 12'hf91: x = 16'h 780; 12'hf92: x = 16'h 777; 12'hf93: x = 16'h 76e; 12'hf94: x = 16'h 765; 12'hf95: x = 16'h 75c; 12'hf96: x = 16'h 753; 12'hf97: x = 16'h 74a; 12'hf98: x = 16'h 741; 12'hf99: x = 16'h 738; 12'hf9a: x = 16'h 72f; 12'hf9b: x = 16'h 726; 12'hf9c: x = 16'h 71d; 12'hf9d: x = 16'h 714; 12'hf9e: x = 16'h 70a; 12'hf9f: x = 16'h 701; 12'hfa0: x = 16'h 6f8; 12'hfa1: x = 16'h 6ee; 12'hfa2: x = 16'h 6e5; 12'hfa3: x = 16'h 6db; 12'hfa4: x = 16'h 6d2; 12'hfa5: x = 16'h 6c8; 12'hfa6: x = 16'h 6be; 12'hfa7: x = 16'h 6b5; 12'hfa8: x = 16'h 6ab; 12'hfa9: x = 16'h 6a1; 12'hfaa: x = 16'h 697; 12'hfab: x = 16'h 68d; 12'hfac: x = 16'h 683; 12'hfad: x = 16'h 679; 12'hfae: x = 16'h 66f; 12'hfaf: x = 16'h 665; 12'hfb0: x = 16'h 65b; 12'hfb1: x = 16'h 650; 12'hfb2: x = 16'h 646; 12'hfb3: x = 16'h 63b; 12'hfb4: x = 16'h 631; 12'hfb5: x = 16'h 626; 12'hfb6: x = 16'h 61c; 12'hfb7: x = 16'h 611; 12'hfb8: x = 16'h 606; 12'hfb9: x = 16'h 5fb; 12'hfba: x = 16'h 5f1; 12'hfbb: x = 16'h 5e6; 12'hfbc: x = 16'h 5da; 12'hfbd: x = 16'h 5cf; 12'hfbe: x = 16'h 5c4; 12'hfbf: x = 16'h 5b9; 12'hfc0: x = 16'h 5ad; 12'hfc1: x = 16'h 5a2; 12'hfc2: x = 16'h 596; 12'hfc3: x = 16'h 58b; 12'hfc4: x = 16'h 57f; 12'hfc5: x = 16'h 573; 12'hfc6: x = 16'h 567; 12'hfc7: x = 16'h 55b; 12'hfc8: x = 16'h 54f; 12'hfc9: x = 16'h 543; 12'hfca: x = 16'h 536; 12'hfcb: x = 16'h 52a; 12'hfcc: x = 16'h 51d; 12'hfcd: x = 16'h 510; 12'hfce: x = 16'h 503; 12'hfcf: x = 16'h 4f6; 12'hfd0: x = 16'h 4e9; 12'hfd1: x = 16'h 4dc; 12'hfd2: x = 16'h 4cf; 12'hfd3: x = 16'h 4c1; 12'hfd4: x = 16'h 4b3; 12'hfd5: x = 16'h 4a6; 12'hfd6: x = 16'h 498; 12'hfd7: x = 16'h 48a; 12'hfd8: x = 16'h 47b; 12'hfd9: x = 16'h 46d; 12'hfda: x = 16'h 45e; 12'hfdb: x = 16'h 44f; 12'hfdc: x = 16'h 440; 12'hfdd: x = 16'h 431; 12'hfde: x = 16'h 421; 12'hfdf: x = 16'h 411; 12'hfe0: x = 16'h 402; 12'hfe1: x = 16'h 3f1; 12'hfe2: x = 16'h 3e1; 12'hfe3: x = 16'h 3d0; 12'hfe4: x = 16'h 3bf; 12'hfe5: x = 16'h 3ae; 12'hfe6: x = 16'h 39c; 12'hfe7: x = 16'h 38a; 12'hfe8: x = 16'h 378; 12'hfe9: x = 16'h 365; 12'hfea: x = 16'h 352; 12'hfeb: x = 16'h 33e; 12'hfec: x = 16'h 32a; 12'hfed: x = 16'h 315; 12'hfee: x = 16'h 300; 12'hfef: x = 16'h 2eb; 12'hff0: x = 16'h 2d4; 12'hff1: x = 16'h 2bd; 12'hff2: x = 16'h 2a5; 12'hff3: x = 16'h 28d; 12'hff4: x = 16'h 273; 12'hff5: x = 16'h 258; 12'hff6: x = 16'h 23c; 12'hff7: x = 16'h 21f; 12'hff8: x = 16'h 200; 12'hff9: x = 16'h 1df; 12'hffa: x = 16'h 1bb; 12'hffb: x = 16'h 194; 12'hffc: x = 16'h 16a; 12'hffd: x = 16'h 139; 12'hffe: x = 16'h 100; 12'hfff: x = 16'h  b5; 
		endcase
	end
endmodule

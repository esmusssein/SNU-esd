module cosin (
	input	[9:0] data_in,
	output [15:0] cos_x_out
);

	reg [15:0] x;
	
	assign cos_x_out = x;
	
	always @(*) begin
		case(data_in)
		10'h  1: x = 16'hffff; 10'h  2: x = 16'hfffe; 10'h  3: x = 16'hfffd; 10'h  4: x = 16'hfffb; 10'h  5: x = 16'hfff8; 10'h  6: x = 16'hfff4; 10'h  7: x = 16'hfff0; 10'h  8: x = 16'hffec; 10'h  9: x = 16'hffe7; 10'h  a: x = 16'hffe1; 10'h  b: x = 16'hffda; 10'h  c: x = 16'hffd3; 10'h  d: x = 16'hffcb; 10'h  e: x = 16'hffc3; 10'h  f: x = 16'hffba; 10'h 10: x = 16'hffb1; 10'h 11: x = 16'hffa6; 10'h 12: x = 16'hff9c; 10'h 13: x = 16'hff90; 10'h 14: x = 16'hff84; 10'h 15: x = 16'hff78; 10'h 16: x = 16'hff6a; 10'h 17: x = 16'hff5c; 10'h 18: x = 16'hff4e; 10'h 19: x = 16'hff3f; 10'h 1a: x = 16'hff2f; 10'h 1b: x = 16'hff1f; 10'h 1c: x = 16'hff0e; 10'h 1d: x = 16'hfefc; 10'h 1e: x = 16'hfeea; 10'h 1f: x = 16'hfed7; 10'h 20: x = 16'hfec4; 10'h 21: x = 16'hfeb0; 10'h 22: x = 16'hfe9b; 10'h 23: x = 16'hfe86; 10'h 24: x = 16'hfe70; 10'h 25: x = 16'hfe5a; 10'h 26: x = 16'hfe43; 10'h 27: x = 16'hfe2b; 10'h 28: x = 16'hfe13; 10'h 29: x = 16'hfdfa; 10'h 2a: x = 16'hfde0; 10'h 2b: x = 16'hfdc6; 10'h 2c: x = 16'hfdab; 10'h 2d: x = 16'hfd90; 10'h 2e: x = 16'hfd74; 10'h 2f: x = 16'hfd57; 10'h 30: x = 16'hfd3a; 10'h 31: x = 16'hfd1c; 10'h 32: x = 16'hfcfe; 10'h 33: x = 16'hfcdf; 10'h 34: x = 16'hfcbf; 10'h 35: x = 16'hfc9f; 10'h 36: x = 16'hfc7e; 10'h 37: x = 16'hfc5d; 10'h 38: x = 16'hfc3b; 10'h 39: x = 16'hfc18; 10'h 3a: x = 16'hfbf5; 10'h 3b: x = 16'hfbd1; 10'h 3c: x = 16'hfbac; 10'h 3d: x = 16'hfb87; 10'h 3e: x = 16'hfb61; 10'h 3f: x = 16'hfb3b; 10'h 40: x = 16'hfb14; 10'h 41: x = 16'hfaed; 10'h 42: x = 16'hfac5; 10'h 43: x = 16'hfa9c; 10'h 44: x = 16'hfa73; 10'h 45: x = 16'hfa49; 10'h 46: x = 16'hfa1e; 10'h 47: x = 16'hf9f3; 10'h 48: x = 16'hf9c7; 10'h 49: x = 16'hf99b; 10'h 4a: x = 16'hf96e; 10'h 4b: x = 16'hf940; 10'h 4c: x = 16'hf912; 10'h 4d: x = 16'hf8e3; 10'h 4e: x = 16'hf8b4; 10'h 4f: x = 16'hf884; 10'h 50: x = 16'hf853; 10'h 51: x = 16'hf822; 10'h 52: x = 16'hf7f1; 10'h 53: x = 16'hf7be; 10'h 54: x = 16'hf78b; 10'h 55: x = 16'hf758; 10'h 56: x = 16'hf724; 10'h 57: x = 16'hf6ef; 10'h 58: x = 16'hf6ba; 10'h 59: x = 16'hf684; 10'h 5a: x = 16'hf64d; 10'h 5b: x = 16'hf616; 10'h 5c: x = 16'hf5de; 10'h 5d: x = 16'hf5a6; 10'h 5e: x = 16'hf56d; 10'h 5f: x = 16'hf534; 10'h 60: x = 16'hf4fa; 10'h 61: x = 16'hf4bf; 10'h 62: x = 16'hf484; 10'h 63: x = 16'hf448; 10'h 64: x = 16'hf40b; 10'h 65: x = 16'hf3ce; 10'h 66: x = 16'hf391; 10'h 67: x = 16'hf353; 10'h 68: x = 16'hf314; 10'h 69: x = 16'hf2d4; 10'h 6a: x = 16'hf294; 10'h 6b: x = 16'hf254; 10'h 6c: x = 16'hf213; 10'h 6d: x = 16'hf1d1; 10'h 6e: x = 16'hf18f; 10'h 6f: x = 16'hf14c; 10'h 70: x = 16'hf109; 10'h 71: x = 16'hf0c5; 10'h 72: x = 16'hf080; 10'h 73: x = 16'hf03b; 10'h 74: x = 16'heff5; 10'h 75: x = 16'hefaf; 10'h 76: x = 16'hef68; 10'h 77: x = 16'hef20; 10'h 78: x = 16'heed8; 10'h 79: x = 16'hee8f; 10'h 7a: x = 16'hee46; 10'h 7b: x = 16'hedfc; 10'h 7c: x = 16'hedb2; 10'h 7d: x = 16'hed67; 10'h 7e: x = 16'hed1c; 10'h 7f: x = 16'hecd0; 10'h 80: x = 16'hec83; 10'h 81: x = 16'hec36; 10'h 82: x = 16'hebe8; 10'h 83: x = 16'heb99; 10'h 84: x = 16'heb4b; 10'h 85: x = 16'heafb; 10'h 86: x = 16'heaab; 10'h 87: x = 16'hea5a; 10'h 88: x = 16'hea09; 10'h 89: x = 16'he9b7; 10'h 8a: x = 16'he965; 10'h 8b: x = 16'he912; 10'h 8c: x = 16'he8bf; 10'h 8d: x = 16'he86b; 10'h 8e: x = 16'he816; 10'h 8f: x = 16'he7c1; 10'h 90: x = 16'he76b; 10'h 91: x = 16'he715; 10'h 92: x = 16'he6be; 10'h 93: x = 16'he667; 10'h 94: x = 16'he60f; 10'h 95: x = 16'he5b7; 10'h 96: x = 16'he55e; 10'h 97: x = 16'he504; 10'h 98: x = 16'he4aa; 10'h 99: x = 16'he44f; 10'h 9a: x = 16'he3f4; 10'h 9b: x = 16'he398; 10'h 9c: x = 16'he33c; 10'h 9d: x = 16'he2df; 10'h 9e: x = 16'he282; 10'h 9f: x = 16'he224; 10'h a0: x = 16'he1c5; 10'h a1: x = 16'he166; 10'h a2: x = 16'he106; 10'h a3: x = 16'he0a6; 10'h a4: x = 16'he046; 10'h a5: x = 16'hdfe4; 10'h a6: x = 16'hdf83; 10'h a7: x = 16'hdf20; 10'h a8: x = 16'hdebe; 10'h a9: x = 16'hde5a; 10'h aa: x = 16'hddf6; 10'h ab: x = 16'hdd92; 10'h ac: x = 16'hdd2d; 10'h ad: x = 16'hdcc7; 10'h ae: x = 16'hdc61; 10'h af: x = 16'hdbfb; 10'h b0: x = 16'hdb94; 10'h b1: x = 16'hdb2c; 10'h b2: x = 16'hdac4; 10'h b3: x = 16'hda5b; 10'h b4: x = 16'hd9f2; 10'h b5: x = 16'hd988; 10'h b6: x = 16'hd91e; 10'h b7: x = 16'hd8b3; 10'h b8: x = 16'hd848; 10'h b9: x = 16'hd7dc; 10'h ba: x = 16'hd770; 10'h bb: x = 16'hd703; 10'h bc: x = 16'hd695; 10'h bd: x = 16'hd627; 10'h be: x = 16'hd5b9; 10'h bf: x = 16'hd54a; 10'h c0: x = 16'hd4db; 10'h c1: x = 16'hd46b; 10'h c2: x = 16'hd3fa; 10'h c3: x = 16'hd389; 10'h c4: x = 16'hd318; 10'h c5: x = 16'hd2a6; 10'h c6: x = 16'hd233; 10'h c7: x = 16'hd1c0; 10'h c8: x = 16'hd14d; 10'h c9: x = 16'hd0d9; 10'h ca: x = 16'hd064; 10'h cb: x = 16'hcfef; 10'h cc: x = 16'hcf7a; 10'h cd: x = 16'hcf04; 10'h ce: x = 16'hce8d; 10'h cf: x = 16'hce16; 10'h d0: x = 16'hcd9f; 10'h d1: x = 16'hcd26; 10'h d2: x = 16'hccae; 10'h d3: x = 16'hcc35; 10'h d4: x = 16'hcbbb; 10'h d5: x = 16'hcb41; 10'h d6: x = 16'hcac7; 10'h d7: x = 16'hca4c; 10'h d8: x = 16'hc9d1; 10'h d9: x = 16'hc955; 10'h da: x = 16'hc8d8; 10'h db: x = 16'hc85b; 10'h dc: x = 16'hc7de; 10'h dd: x = 16'hc760; 10'h de: x = 16'hc6e2; 10'h df: x = 16'hc663; 10'h e0: x = 16'hc5e4; 10'h e1: x = 16'hc564; 10'h e2: x = 16'hc4e3; 10'h e3: x = 16'hc463; 10'h e4: x = 16'hc3e2; 10'h e5: x = 16'hc360; 10'h e6: x = 16'hc2de; 10'h e7: x = 16'hc25b; 10'h e8: x = 16'hc1d8; 10'h e9: x = 16'hc154; 10'h ea: x = 16'hc0d0; 10'h eb: x = 16'hc04c; 10'h ec: x = 16'hbfc7; 10'h ed: x = 16'hbf41; 10'h ee: x = 16'hbebc; 10'h ef: x = 16'hbe35; 10'h f0: x = 16'hbdae; 10'h f1: x = 16'hbd27; 10'h f2: x = 16'hbca0; 10'h f3: x = 16'hbc17; 10'h f4: x = 16'hbb8f; 10'h f5: x = 16'hbb06; 10'h f6: x = 16'hba7c; 10'h f7: x = 16'hb9f2; 10'h f8: x = 16'hb968; 10'h f9: x = 16'hb8dd; 10'h fa: x = 16'hb852; 10'h fb: x = 16'hb7c6; 10'h fc: x = 16'hb73a; 10'h fd: x = 16'hb6ad; 10'h fe: x = 16'hb620; 10'h ff: x = 16'hb592; 10'h100: x = 16'hb504; 10'h101: x = 16'hb476; 10'h102: x = 16'hb3e7; 10'h103: x = 16'hb358; 10'h104: x = 16'hb2c8; 10'h105: x = 16'hb238; 10'h106: x = 16'hb1a8; 10'h107: x = 16'hb117; 10'h108: x = 16'hb085; 10'h109: x = 16'haff3; 10'h10a: x = 16'haf61; 10'h10b: x = 16'haece; 10'h10c: x = 16'hae3b; 10'h10d: x = 16'hada8; 10'h10e: x = 16'had14; 10'h10f: x = 16'hac80; 10'h110: x = 16'habeb; 10'h111: x = 16'hab56; 10'h112: x = 16'haac0; 10'h113: x = 16'haa2a; 10'h114: x = 16'ha994; 10'h115: x = 16'ha8fd; 10'h116: x = 16'ha866; 10'h117: x = 16'ha7ce; 10'h118: x = 16'ha736; 10'h119: x = 16'ha69d; 10'h11a: x = 16'ha605; 10'h11b: x = 16'ha56b; 10'h11c: x = 16'ha4d2; 10'h11d: x = 16'ha438; 10'h11e: x = 16'ha39d; 10'h11f: x = 16'ha302; 10'h120: x = 16'ha267; 10'h121: x = 16'ha1cb; 10'h122: x = 16'ha12f; 10'h123: x = 16'ha093; 10'h124: x = 16'h9ff6; 10'h125: x = 16'h9f59; 10'h126: x = 16'h9ebc; 10'h127: x = 16'h9e1e; 10'h128: x = 16'h9d7f; 10'h129: x = 16'h9ce1; 10'h12a: x = 16'h9c42; 10'h12b: x = 16'h9ba2; 10'h12c: x = 16'h9b02; 10'h12d: x = 16'h9a62; 10'h12e: x = 16'h99c2; 10'h12f: x = 16'h9921; 10'h130: x = 16'h987f; 10'h131: x = 16'h97de; 10'h132: x = 16'h973c; 10'h133: x = 16'h9699; 10'h134: x = 16'h95f6; 10'h135: x = 16'h9553; 10'h136: x = 16'h94b0; 10'h137: x = 16'h940c; 10'h138: x = 16'h9368; 10'h139: x = 16'h92c3; 10'h13a: x = 16'h921e; 10'h13b: x = 16'h9179; 10'h13c: x = 16'h90d3; 10'h13d: x = 16'h902d; 10'h13e: x = 16'h8f87; 10'h13f: x = 16'h8ee0; 10'h140: x = 16'h8e39; 10'h141: x = 16'h8d92; 10'h142: x = 16'h8cea; 10'h143: x = 16'h8c42; 10'h144: x = 16'h8b9a; 10'h145: x = 16'h8af1; 10'h146: x = 16'h8a48; 10'h147: x = 16'h899f; 10'h148: x = 16'h88f5; 10'h149: x = 16'h884b; 10'h14a: x = 16'h87a1; 10'h14b: x = 16'h86f6; 10'h14c: x = 16'h864b; 10'h14d: x = 16'h85a0; 10'h14e: x = 16'h84f4; 10'h14f: x = 16'h8448; 10'h150: x = 16'h839c; 10'h151: x = 16'h82ef; 10'h152: x = 16'h8242; 10'h153: x = 16'h8195; 10'h154: x = 16'h80e7; 10'h155: x = 16'h803a; 10'h156: x = 16'h7f8b; 10'h157: x = 16'h7edd; 10'h158: x = 16'h7e2e; 10'h159: x = 16'h7d7f; 10'h15a: x = 16'h7cd0; 10'h15b: x = 16'h7c20; 10'h15c: x = 16'h7b70; 10'h15d: x = 16'h7ac0; 10'h15e: x = 16'h7a0f; 10'h15f: x = 16'h795e; 10'h160: x = 16'h78ad; 10'h161: x = 16'h77fb; 10'h162: x = 16'h774a; 10'h163: x = 16'h7698; 10'h164: x = 16'h75e5; 10'h165: x = 16'h7533; 10'h166: x = 16'h7480; 10'h167: x = 16'h73cd; 10'h168: x = 16'h7319; 10'h169: x = 16'h7265; 10'h16a: x = 16'h71b1; 10'h16b: x = 16'h70fd; 10'h16c: x = 16'h7049; 10'h16d: x = 16'h6f94; 10'h16e: x = 16'h6edf; 10'h16f: x = 16'h6e29; 10'h170: x = 16'h6d74; 10'h171: x = 16'h6cbe; 10'h172: x = 16'h6c08; 10'h173: x = 16'h6b51; 10'h174: x = 16'h6a9b; 10'h175: x = 16'h69e4; 10'h176: x = 16'h692d; 10'h177: x = 16'h6875; 10'h178: x = 16'h67bd; 10'h179: x = 16'h6705; 10'h17a: x = 16'h664d; 10'h17b: x = 16'h6595; 10'h17c: x = 16'h64dc; 10'h17d: x = 16'h6423; 10'h17e: x = 16'h636a; 10'h17f: x = 16'h62b1; 10'h180: x = 16'h61f7; 10'h181: x = 16'h613d; 10'h182: x = 16'h6083; 10'h183: x = 16'h5fc9; 10'h184: x = 16'h5f0e; 10'h185: x = 16'h5e53; 10'h186: x = 16'h5d98; 10'h187: x = 16'h5cdd; 10'h188: x = 16'h5c22; 10'h189: x = 16'h5b66; 10'h18a: x = 16'h5aaa; 10'h18b: x = 16'h59ee; 10'h18c: x = 16'h5931; 10'h18d: x = 16'h5875; 10'h18e: x = 16'h57b8; 10'h18f: x = 16'h56fb; 10'h190: x = 16'h563e; 10'h191: x = 16'h5581; 10'h192: x = 16'h54c3; 10'h193: x = 16'h5405; 10'h194: x = 16'h5347; 10'h195: x = 16'h5289; 10'h196: x = 16'h51ca; 10'h197: x = 16'h510c; 10'h198: x = 16'h504d; 10'h199: x = 16'h4f8e; 10'h19a: x = 16'h4ecf; 10'h19b: x = 16'h4e0f; 10'h19c: x = 16'h4d50; 10'h19d: x = 16'h4c90; 10'h19e: x = 16'h4bd0; 10'h19f: x = 16'h4b10; 10'h1a0: x = 16'h4a50; 10'h1a1: x = 16'h498f; 10'h1a2: x = 16'h48ce; 10'h1a3: x = 16'h480e; 10'h1a4: x = 16'h474d; 10'h1a5: x = 16'h468b; 10'h1a6: x = 16'h45ca; 10'h1a7: x = 16'h4508; 10'h1a8: x = 16'h4447; 10'h1a9: x = 16'h4385; 10'h1aa: x = 16'h42c3; 10'h1ab: x = 16'h4201; 10'h1ac: x = 16'h413e; 10'h1ad: x = 16'h407c; 10'h1ae: x = 16'h3fb9; 10'h1af: x = 16'h3ef6; 10'h1b0: x = 16'h3e33; 10'h1b1: x = 16'h3d70; 10'h1b2: x = 16'h3cad; 10'h1b3: x = 16'h3bea; 10'h1b4: x = 16'h3b26; 10'h1b5: x = 16'h3a62; 10'h1b6: x = 16'h399f; 10'h1b7: x = 16'h38db; 10'h1b8: x = 16'h3817; 10'h1b9: x = 16'h3752; 10'h1ba: x = 16'h368e; 10'h1bb: x = 16'h35c9; 10'h1bc: x = 16'h3505; 10'h1bd: x = 16'h3440; 10'h1be: x = 16'h337b; 10'h1bf: x = 16'h32b6; 10'h1c0: x = 16'h31f1; 10'h1c1: x = 16'h312c; 10'h1c2: x = 16'h3066; 10'h1c3: x = 16'h2fa1; 10'h1c4: x = 16'h2edb; 10'h1c5: x = 16'h2e15; 10'h1c6: x = 16'h2d50; 10'h1c7: x = 16'h2c8a; 10'h1c8: x = 16'h2bc4; 10'h1c9: x = 16'h2afe; 10'h1ca: x = 16'h2a37; 10'h1cb: x = 16'h2971; 10'h1cc: x = 16'h28aa; 10'h1cd: x = 16'h27e4; 10'h1ce: x = 16'h271d; 10'h1cf: x = 16'h2656; 10'h1d0: x = 16'h2590; 10'h1d1: x = 16'h24c9; 10'h1d2: x = 16'h2402; 10'h1d3: x = 16'h233b; 10'h1d4: x = 16'h2273; 10'h1d5: x = 16'h21ac; 10'h1d6: x = 16'h20e5; 10'h1d7: x = 16'h201d; 10'h1d8: x = 16'h1f56; 10'h1d9: x = 16'h1e8e; 10'h1da: x = 16'h1dc7; 10'h1db: x = 16'h1cff; 10'h1dc: x = 16'h1c37; 10'h1dd: x = 16'h1b6f; 10'h1de: x = 16'h1aa7; 10'h1df: x = 16'h19df; 10'h1e0: x = 16'h1917; 10'h1e1: x = 16'h184f; 10'h1e2: x = 16'h1787; 10'h1e3: x = 16'h16bf; 10'h1e4: x = 16'h15f6; 10'h1e5: x = 16'h152e; 10'h1e6: x = 16'h1466; 10'h1e7: x = 16'h139d; 10'h1e8: x = 16'h12d5; 10'h1e9: x = 16'h120c; 10'h1ea: x = 16'h1144; 10'h1eb: x = 16'h107b; 10'h1ec: x = 16'h fb2; 10'h1ed: x = 16'h eea; 10'h1ee: x = 16'h e21; 10'h1ef: x = 16'h d58; 10'h1f0: x = 16'h c8f; 10'h1f1: x = 16'h bc6; 10'h1f2: x = 16'h afe; 10'h1f3: x = 16'h a35; 10'h1f4: x = 16'h 96c; 10'h1f5: x = 16'h 8a3; 10'h1f6: x = 16'h 7da; 10'h1f7: x = 16'h 711; 10'h1f8: x = 16'h 648; 10'h1f9: x = 16'h 57f; 10'h1fa: x = 16'h 4b6; 10'h1fb: x = 16'h 3ed; 10'h1fc: x = 16'h 324; 10'h1fd: x = 16'h 25b; 10'h1fe: x = 16'h 192; 10'h1ff: x = 16'h  c9; 10'h200: x = 16'h   0; 10'h201: x = 16'hffffff37; 10'h202: x = 16'hfffffe6e; 10'h203: x = 16'hfffffda5; 10'h204: x = 16'hfffffcdc; 10'h205: x = 16'hfffffc13; 10'h206: x = 16'hfffffb4a; 10'h207: x = 16'hfffffa81; 10'h208: x = 16'hfffff9b8; 10'h209: x = 16'hfffff8ef; 10'h20a: x = 16'hfffff826; 10'h20b: x = 16'hfffff75d; 10'h20c: x = 16'hfffff694; 10'h20d: x = 16'hfffff5cb; 10'h20e: x = 16'hfffff502; 10'h20f: x = 16'hfffff43a; 10'h210: x = 16'hfffff371; 10'h211: x = 16'hfffff2a8; 10'h212: x = 16'hfffff1df; 10'h213: x = 16'hfffff116; 10'h214: x = 16'hfffff04e; 10'h215: x = 16'hffffef85; 10'h216: x = 16'hffffeebc; 10'h217: x = 16'hffffedf4; 10'h218: x = 16'hffffed2b; 10'h219: x = 16'hffffec63; 10'h21a: x = 16'hffffeb9a; 10'h21b: x = 16'hffffead2; 10'h21c: x = 16'hffffea0a; 10'h21d: x = 16'hffffe941; 10'h21e: x = 16'hffffe879; 10'h21f: x = 16'hffffe7b1; 10'h220: x = 16'hffffe6e9; 10'h221: x = 16'hffffe621; 10'h222: x = 16'hffffe559; 10'h223: x = 16'hffffe491; 10'h224: x = 16'hffffe3c9; 10'h225: x = 16'hffffe301; 10'h226: x = 16'hffffe239; 10'h227: x = 16'hffffe172; 10'h228: x = 16'hffffe0aa; 10'h229: x = 16'hffffdfe3; 10'h22a: x = 16'hffffdf1b; 10'h22b: x = 16'hffffde54; 10'h22c: x = 16'hffffdd8d; 10'h22d: x = 16'hffffdcc5; 10'h22e: x = 16'hffffdbfe; 10'h22f: x = 16'hffffdb37; 10'h230: x = 16'hffffda70; 10'h231: x = 16'hffffd9aa; 10'h232: x = 16'hffffd8e3; 10'h233: x = 16'hffffd81c; 10'h234: x = 16'hffffd756; 10'h235: x = 16'hffffd68f; 10'h236: x = 16'hffffd5c9; 10'h237: x = 16'hffffd502; 10'h238: x = 16'hffffd43c; 10'h239: x = 16'hffffd376; 10'h23a: x = 16'hffffd2b0; 10'h23b: x = 16'hffffd1eb; 10'h23c: x = 16'hffffd125; 10'h23d: x = 16'hffffd05f; 10'h23e: x = 16'hffffcf9a; 10'h23f: x = 16'hffffced4; 10'h240: x = 16'hffffce0f; 10'h241: x = 16'hffffcd4a; 10'h242: x = 16'hffffcc85; 10'h243: x = 16'hffffcbc0; 10'h244: x = 16'hffffcafb; 10'h245: x = 16'hffffca37; 10'h246: x = 16'hffffc972; 10'h247: x = 16'hffffc8ae; 10'h248: x = 16'hffffc7e9; 10'h249: x = 16'hffffc725; 10'h24a: x = 16'hffffc661; 10'h24b: x = 16'hffffc59e; 10'h24c: x = 16'hffffc4da; 10'h24d: x = 16'hffffc416; 10'h24e: x = 16'hffffc353; 10'h24f: x = 16'hffffc290; 10'h250: x = 16'hffffc1cd; 10'h251: x = 16'hffffc10a; 10'h252: x = 16'hffffc047; 10'h253: x = 16'hffffbf84; 10'h254: x = 16'hffffbec2; 10'h255: x = 16'hffffbdff; 10'h256: x = 16'hffffbd3d; 10'h257: x = 16'hffffbc7b; 10'h258: x = 16'hffffbbb9; 10'h259: x = 16'hffffbaf8; 10'h25a: x = 16'hffffba36; 10'h25b: x = 16'hffffb975; 10'h25c: x = 16'hffffb8b3; 10'h25d: x = 16'hffffb7f2; 10'h25e: x = 16'hffffb732; 10'h25f: x = 16'hffffb671; 10'h260: x = 16'hffffb5b0; 10'h261: x = 16'hffffb4f0; 10'h262: x = 16'hffffb430; 10'h263: x = 16'hffffb370; 10'h264: x = 16'hffffb2b0; 10'h265: x = 16'hffffb1f1; 10'h266: x = 16'hffffb131; 10'h267: x = 16'hffffb072; 10'h268: x = 16'hffffafb3; 10'h269: x = 16'hffffaef4; 10'h26a: x = 16'hffffae36; 10'h26b: x = 16'hffffad77; 10'h26c: x = 16'hffffacb9; 10'h26d: x = 16'hffffabfb; 10'h26e: x = 16'hffffab3d; 10'h26f: x = 16'hffffaa7f; 10'h270: x = 16'hffffa9c2; 10'h271: x = 16'hffffa905; 10'h272: x = 16'hffffa848; 10'h273: x = 16'hffffa78b; 10'h274: x = 16'hffffa6cf; 10'h275: x = 16'hffffa612; 10'h276: x = 16'hffffa556; 10'h277: x = 16'hffffa49a; 10'h278: x = 16'hffffa3de; 10'h279: x = 16'hffffa323; 10'h27a: x = 16'hffffa268; 10'h27b: x = 16'hffffa1ad; 10'h27c: x = 16'hffffa0f2; 10'h27d: x = 16'hffffa037; 10'h27e: x = 16'hffff9f7d; 10'h27f: x = 16'hffff9ec3; 10'h280: x = 16'hffff9e09; 10'h281: x = 16'hffff9d4f; 10'h282: x = 16'hffff9c96; 10'h283: x = 16'hffff9bdd; 10'h284: x = 16'hffff9b24; 10'h285: x = 16'hffff9a6b; 10'h286: x = 16'hffff99b3; 10'h287: x = 16'hffff98fb; 10'h288: x = 16'hffff9843; 10'h289: x = 16'hffff978b; 10'h28a: x = 16'hffff96d3; 10'h28b: x = 16'hffff961c; 10'h28c: x = 16'hffff9565; 10'h28d: x = 16'hffff94af; 10'h28e: x = 16'hffff93f8; 10'h28f: x = 16'hffff9342; 10'h290: x = 16'hffff928c; 10'h291: x = 16'hffff91d7; 10'h292: x = 16'hffff9121; 10'h293: x = 16'hffff906c; 10'h294: x = 16'hffff8fb7; 10'h295: x = 16'hffff8f03; 10'h296: x = 16'hffff8e4f; 10'h297: x = 16'hffff8d9b; 10'h298: x = 16'hffff8ce7; 10'h299: x = 16'hffff8c33; 10'h29a: x = 16'hffff8b80; 10'h29b: x = 16'hffff8acd; 10'h29c: x = 16'hffff8a1b; 10'h29d: x = 16'hffff8968; 10'h29e: x = 16'hffff88b6; 10'h29f: x = 16'hffff8805; 10'h2a0: x = 16'hffff8753; 10'h2a1: x = 16'hffff86a2; 10'h2a2: x = 16'hffff85f1; 10'h2a3: x = 16'hffff8540; 10'h2a4: x = 16'hffff8490; 10'h2a5: x = 16'hffff83e0; 10'h2a6: x = 16'hffff8330; 10'h2a7: x = 16'hffff8281; 10'h2a8: x = 16'hffff81d2; 10'h2a9: x = 16'hffff8123; 10'h2aa: x = 16'hffff8075; 10'h2ab: x = 16'hffff7fc6; 10'h2ac: x = 16'hffff7f19; 10'h2ad: x = 16'hffff7e6b; 10'h2ae: x = 16'hffff7dbe; 10'h2af: x = 16'hffff7d11; 10'h2b0: x = 16'hffff7c64; 10'h2b1: x = 16'hffff7bb8; 10'h2b2: x = 16'hffff7b0c; 10'h2b3: x = 16'hffff7a60; 10'h2b4: x = 16'hffff79b5; 10'h2b5: x = 16'hffff790a; 10'h2b6: x = 16'hffff785f; 10'h2b7: x = 16'hffff77b5; 10'h2b8: x = 16'hffff770b; 10'h2b9: x = 16'hffff7661; 10'h2ba: x = 16'hffff75b8; 10'h2bb: x = 16'hffff750f; 10'h2bc: x = 16'hffff7466; 10'h2bd: x = 16'hffff73be; 10'h2be: x = 16'hffff7316; 10'h2bf: x = 16'hffff726e; 10'h2c0: x = 16'hffff71c7; 10'h2c1: x = 16'hffff7120; 10'h2c2: x = 16'hffff7079; 10'h2c3: x = 16'hffff6fd3; 10'h2c4: x = 16'hffff6f2d; 10'h2c5: x = 16'hffff6e87; 10'h2c6: x = 16'hffff6de2; 10'h2c7: x = 16'hffff6d3d; 10'h2c8: x = 16'hffff6c98; 10'h2c9: x = 16'hffff6bf4; 10'h2ca: x = 16'hffff6b50; 10'h2cb: x = 16'hffff6aad; 10'h2cc: x = 16'hffff6a0a; 10'h2cd: x = 16'hffff6967; 10'h2ce: x = 16'hffff68c4; 10'h2cf: x = 16'hffff6822; 10'h2d0: x = 16'hffff6781; 10'h2d1: x = 16'hffff66df; 10'h2d2: x = 16'hffff663e; 10'h2d3: x = 16'hffff659e; 10'h2d4: x = 16'hffff64fe; 10'h2d5: x = 16'hffff645e; 10'h2d6: x = 16'hffff63be; 10'h2d7: x = 16'hffff631f; 10'h2d8: x = 16'hffff6281; 10'h2d9: x = 16'hffff61e2; 10'h2da: x = 16'hffff6144; 10'h2db: x = 16'hffff60a7; 10'h2dc: x = 16'hffff600a; 10'h2dd: x = 16'hffff5f6d; 10'h2de: x = 16'hffff5ed1; 10'h2df: x = 16'hffff5e35; 10'h2e0: x = 16'hffff5d99; 10'h2e1: x = 16'hffff5cfe; 10'h2e2: x = 16'hffff5c63; 10'h2e3: x = 16'hffff5bc8; 10'h2e4: x = 16'hffff5b2e; 10'h2e5: x = 16'hffff5a95; 10'h2e6: x = 16'hffff59fb; 10'h2e7: x = 16'hffff5963; 10'h2e8: x = 16'hffff58ca; 10'h2e9: x = 16'hffff5832; 10'h2ea: x = 16'hffff579a; 10'h2eb: x = 16'hffff5703; 10'h2ec: x = 16'hffff566c; 10'h2ed: x = 16'hffff55d6; 10'h2ee: x = 16'hffff5540; 10'h2ef: x = 16'hffff54aa; 10'h2f0: x = 16'hffff5415; 10'h2f1: x = 16'hffff5380; 10'h2f2: x = 16'hffff52ec; 10'h2f3: x = 16'hffff5258; 10'h2f4: x = 16'hffff51c5; 10'h2f5: x = 16'hffff5132; 10'h2f6: x = 16'hffff509f; 10'h2f7: x = 16'hffff500d; 10'h2f8: x = 16'hffff4f7b; 10'h2f9: x = 16'hffff4ee9; 10'h2fa: x = 16'hffff4e58; 10'h2fb: x = 16'hffff4dc8; 10'h2fc: x = 16'hffff4d38; 10'h2fd: x = 16'hffff4ca8; 10'h2fe: x = 16'hffff4c19; 10'h2ff: x = 16'hffff4b8a; 10'h300: x = 16'hffff4afc; 10'h301: x = 16'hffff4a6e; 10'h302: x = 16'hffff49e0; 10'h303: x = 16'hffff4953; 10'h304: x = 16'hffff48c6; 10'h305: x = 16'hffff483a; 10'h306: x = 16'hffff47ae; 10'h307: x = 16'hffff4723; 10'h308: x = 16'hffff4698; 10'h309: x = 16'hffff460e; 10'h30a: x = 16'hffff4584; 10'h30b: x = 16'hffff44fa; 10'h30c: x = 16'hffff4471; 10'h30d: x = 16'hffff43e9; 10'h30e: x = 16'hffff4360; 10'h30f: x = 16'hffff42d9; 10'h310: x = 16'hffff4252; 10'h311: x = 16'hffff41cb; 10'h312: x = 16'hffff4144; 10'h313: x = 16'hffff40bf; 10'h314: x = 16'hffff4039; 10'h315: x = 16'hffff3fb4; 10'h316: x = 16'hffff3f30; 10'h317: x = 16'hffff3eac; 10'h318: x = 16'hffff3e28; 10'h319: x = 16'hffff3da5; 10'h31a: x = 16'hffff3d22; 10'h31b: x = 16'hffff3ca0; 10'h31c: x = 16'hffff3c1e; 10'h31d: x = 16'hffff3b9d; 10'h31e: x = 16'hffff3b1d; 10'h31f: x = 16'hffff3a9c; 10'h320: x = 16'hffff3a1c; 10'h321: x = 16'hffff399d; 10'h322: x = 16'hffff391e; 10'h323: x = 16'hffff38a0; 10'h324: x = 16'hffff3822; 10'h325: x = 16'hffff37a5; 10'h326: x = 16'hffff3728; 10'h327: x = 16'hffff36ab; 10'h328: x = 16'hffff362f; 10'h329: x = 16'hffff35b4; 10'h32a: x = 16'hffff3539; 10'h32b: x = 16'hffff34bf; 10'h32c: x = 16'hffff3445; 10'h32d: x = 16'hffff33cb; 10'h32e: x = 16'hffff3352; 10'h32f: x = 16'hffff32da; 10'h330: x = 16'hffff3261; 10'h331: x = 16'hffff31ea; 10'h332: x = 16'hffff3173; 10'h333: x = 16'hffff30fc; 10'h334: x = 16'hffff3086; 10'h335: x = 16'hffff3011; 10'h336: x = 16'hffff2f9c; 10'h337: x = 16'hffff2f27; 10'h338: x = 16'hffff2eb3; 10'h339: x = 16'hffff2e40; 10'h33a: x = 16'hffff2dcd; 10'h33b: x = 16'hffff2d5a; 10'h33c: x = 16'hffff2ce8; 10'h33d: x = 16'hffff2c77; 10'h33e: x = 16'hffff2c06; 10'h33f: x = 16'hffff2b95; 10'h340: x = 16'hffff2b25; 10'h341: x = 16'hffff2ab6; 10'h342: x = 16'hffff2a47; 10'h343: x = 16'hffff29d9; 10'h344: x = 16'hffff296b; 10'h345: x = 16'hffff28fd; 10'h346: x = 16'hffff2890; 10'h347: x = 16'hffff2824; 10'h348: x = 16'hffff27b8; 10'h349: x = 16'hffff274d; 10'h34a: x = 16'hffff26e2; 10'h34b: x = 16'hffff2678; 10'h34c: x = 16'hffff260e; 10'h34d: x = 16'hffff25a5; 10'h34e: x = 16'hffff253c; 10'h34f: x = 16'hffff24d4; 10'h350: x = 16'hffff246c; 10'h351: x = 16'hffff2405; 10'h352: x = 16'hffff239f; 10'h353: x = 16'hffff2339; 10'h354: x = 16'hffff22d3; 10'h355: x = 16'hffff226e; 10'h356: x = 16'hffff220a; 10'h357: x = 16'hffff21a6; 10'h358: x = 16'hffff2142; 10'h359: x = 16'hffff20e0; 10'h35a: x = 16'hffff207d; 10'h35b: x = 16'hffff201c; 10'h35c: x = 16'hffff1fba; 10'h35d: x = 16'hffff1f5a; 10'h35e: x = 16'hffff1efa; 10'h35f: x = 16'hffff1e9a; 10'h360: x = 16'hffff1e3b; 10'h361: x = 16'hffff1ddc; 10'h362: x = 16'hffff1d7e; 10'h363: x = 16'hffff1d21; 10'h364: x = 16'hffff1cc4; 10'h365: x = 16'hffff1c68; 10'h366: x = 16'hffff1c0c; 10'h367: x = 16'hffff1bb1; 10'h368: x = 16'hffff1b56; 10'h369: x = 16'hffff1afc; 10'h36a: x = 16'hffff1aa2; 10'h36b: x = 16'hffff1a49; 10'h36c: x = 16'hffff19f1; 10'h36d: x = 16'hffff1999; 10'h36e: x = 16'hffff1942; 10'h36f: x = 16'hffff18eb; 10'h370: x = 16'hffff1895; 10'h371: x = 16'hffff183f; 10'h372: x = 16'hffff17ea; 10'h373: x = 16'hffff1795; 10'h374: x = 16'hffff1741; 10'h375: x = 16'hffff16ee; 10'h376: x = 16'hffff169b; 10'h377: x = 16'hffff1649; 10'h378: x = 16'hffff15f7; 10'h379: x = 16'hffff15a6; 10'h37a: x = 16'hffff1555; 10'h37b: x = 16'hffff1505; 10'h37c: x = 16'hffff14b5; 10'h37d: x = 16'hffff1467; 10'h37e: x = 16'hffff1418; 10'h37f: x = 16'hffff13ca; 10'h380: x = 16'hffff137d; 10'h381: x = 16'hffff1330; 10'h382: x = 16'hffff12e4; 10'h383: x = 16'hffff1299; 10'h384: x = 16'hffff124e; 10'h385: x = 16'hffff1204; 10'h386: x = 16'hffff11ba; 10'h387: x = 16'hffff1171; 10'h388: x = 16'hffff1128; 10'h389: x = 16'hffff10e0; 10'h38a: x = 16'hffff1098; 10'h38b: x = 16'hffff1051; 10'h38c: x = 16'hffff100b; 10'h38d: x = 16'hffff0fc5; 10'h38e: x = 16'hffff0f80; 10'h38f: x = 16'hffff0f3b; 10'h390: x = 16'hffff0ef7; 10'h391: x = 16'hffff0eb4; 10'h392: x = 16'hffff0e71; 10'h393: x = 16'hffff0e2f; 10'h394: x = 16'hffff0ded; 10'h395: x = 16'hffff0dac; 10'h396: x = 16'hffff0d6c; 10'h397: x = 16'hffff0d2c; 10'h398: x = 16'hffff0cec; 10'h399: x = 16'hffff0cad; 10'h39a: x = 16'hffff0c6f; 10'h39b: x = 16'hffff0c32; 10'h39c: x = 16'hffff0bf5; 10'h39d: x = 16'hffff0bb8; 10'h39e: x = 16'hffff0b7c; 10'h39f: x = 16'hffff0b41; 10'h3a0: x = 16'hffff0b06; 10'h3a1: x = 16'hffff0acc; 10'h3a2: x = 16'hffff0a93; 10'h3a3: x = 16'hffff0a5a; 10'h3a4: x = 16'hffff0a22; 10'h3a5: x = 16'hffff09ea; 10'h3a6: x = 16'hffff09b3; 10'h3a7: x = 16'hffff097c; 10'h3a8: x = 16'hffff0946; 10'h3a9: x = 16'hffff0911; 10'h3aa: x = 16'hffff08dc; 10'h3ab: x = 16'hffff08a8; 10'h3ac: x = 16'hffff0875; 10'h3ad: x = 16'hffff0842; 10'h3ae: x = 16'hffff080f; 10'h3af: x = 16'hffff07de; 10'h3b0: x = 16'hffff07ad; 10'h3b1: x = 16'hffff077c; 10'h3b2: x = 16'hffff074c; 10'h3b3: x = 16'hffff071d; 10'h3b4: x = 16'hffff06ee; 10'h3b5: x = 16'hffff06c0; 10'h3b6: x = 16'hffff0692; 10'h3b7: x = 16'hffff0665; 10'h3b8: x = 16'hffff0639; 10'h3b9: x = 16'hffff060d; 10'h3ba: x = 16'hffff05e2; 10'h3bb: x = 16'hffff05b7; 10'h3bc: x = 16'hffff058d; 10'h3bd: x = 16'hffff0564; 10'h3be: x = 16'hffff053b; 10'h3bf: x = 16'hffff0513; 10'h3c0: x = 16'hffff04ec; 10'h3c1: x = 16'hffff04c5; 10'h3c2: x = 16'hffff049f; 10'h3c3: x = 16'hffff0479; 10'h3c4: x = 16'hffff0454; 10'h3c5: x = 16'hffff042f; 10'h3c6: x = 16'hffff040b; 10'h3c7: x = 16'hffff03e8; 10'h3c8: x = 16'hffff03c5; 10'h3c9: x = 16'hffff03a3; 10'h3ca: x = 16'hffff0382; 10'h3cb: x = 16'hffff0361; 10'h3cc: x = 16'hffff0341; 10'h3cd: x = 16'hffff0321; 10'h3ce: x = 16'hffff0302; 10'h3cf: x = 16'hffff02e4; 10'h3d0: x = 16'hffff02c6; 10'h3d1: x = 16'hffff02a9; 10'h3d2: x = 16'hffff028c; 10'h3d3: x = 16'hffff0270; 10'h3d4: x = 16'hffff0255; 10'h3d5: x = 16'hffff023a; 10'h3d6: x = 16'hffff0220; 10'h3d7: x = 16'hffff0206; 10'h3d8: x = 16'hffff01ed; 10'h3d9: x = 16'hffff01d5; 10'h3da: x = 16'hffff01bd; 10'h3db: x = 16'hffff01a6; 10'h3dc: x = 16'hffff0190; 10'h3dd: x = 16'hffff017a; 10'h3de: x = 16'hffff0165; 10'h3df: x = 16'hffff0150; 10'h3e0: x = 16'hffff013c; 10'h3e1: x = 16'hffff0129; 10'h3e2: x = 16'hffff0116; 10'h3e3: x = 16'hffff0104; 10'h3e4: x = 16'hffff00f2; 10'h3e5: x = 16'hffff00e1; 10'h3e6: x = 16'hffff00d1; 10'h3e7: x = 16'hffff00c1; 10'h3e8: x = 16'hffff00b2; 10'h3e9: x = 16'hffff00a4; 10'h3ea: x = 16'hffff0096; 10'h3eb: x = 16'hffff0088; 10'h3ec: x = 16'hffff007c; 10'h3ed: x = 16'hffff0070; 10'h3ee: x = 16'hffff0064; 10'h3ef: x = 16'hffff005a; 10'h3f0: x = 16'hffff004f; 10'h3f1: x = 16'hffff0046; 10'h3f2: x = 16'hffff003d; 10'h3f3: x = 16'hffff0035; 10'h3f4: x = 16'hffff002d; 10'h3f5: x = 16'hffff0026; 10'h3f6: x = 16'hffff001f; 10'h3f7: x = 16'hffff0019; 10'h3f8: x = 16'hffff0014; 10'h3f9: x = 16'hffff0010; 10'h3fa: x = 16'hffff000c; 10'h3fb: x = 16'hffff0008; 10'h3fc: x = 16'hffff0005; 10'h3fd: x = 16'hffff0003; 10'h3fe: x = 16'hffff0002; 10'h3ff: x = 16'hffff0001; 			
		default: x = 16'h0000;
		endcase
	end
endmodule

module sqrt_log (
	input	[13:0] data_in,
	output [15:0] data_out
);
	reg [15:0] x;
	
	assign data_out = x;
	
	always @(*) begin
		case(data_in)
		14'h   1: x = 16'h8cf9; 14'h   2: x = 16'h87d8; 14'h   3: x = 16'h84c1; 14'h   4: x = 16'h8284; 14'h   5: x = 16'h80c1; 14'h   6: x = 16'h7f4b; 14'h   7: x = 16'h7e0c; 14'h   8: x = 16'h7cf5; 14'h   9: x = 16'h7bfd; 14'h   a: x = 16'h7b1e; 14'h   b: x = 16'h7a52; 14'h   c: x = 16'h7997; 14'h   d: x = 16'h78ea; 14'h   e: x = 16'h7849; 14'h   f: x = 16'h77b2; 14'h  10: x = 16'h7725; 14'h  11: x = 16'h769f; 14'h  12: x = 16'h7620; 14'h  13: x = 16'h75a8; 14'h  14: x = 16'h7536; 14'h  15: x = 16'h74c8; 14'h  16: x = 16'h7460; 14'h  17: x = 16'h73fc; 14'h  18: x = 16'h739b; 14'h  19: x = 16'h733e; 14'h  1a: x = 16'h72e5; 14'h  1b: x = 16'h728f; 14'h  1c: x = 16'h723c; 14'h  1d: x = 16'h71eb; 14'h  1e: x = 16'h719d; 14'h  1f: x = 16'h7151; 14'h  20: x = 16'h7108; 14'h  21: x = 16'h70c0; 14'h  22: x = 16'h707b; 14'h  23: x = 16'h7037; 14'h  24: x = 16'h6ff5; 14'h  25: x = 16'h6fb5; 14'h  26: x = 16'h6f76; 14'h  27: x = 16'h6f39; 14'h  28: x = 16'h6efd; 14'h  29: x = 16'h6ec3; 14'h  2a: x = 16'h6e8a; 14'h  2b: x = 16'h6e52; 14'h  2c: x = 16'h6e1b; 14'h  2d: x = 16'h6de6; 14'h  2e: x = 16'h6db1; 14'h  2f: x = 16'h6d7e; 14'h  30: x = 16'h6d4b; 14'h  31: x = 16'h6d1a; 14'h  32: x = 16'h6ce9; 14'h  33: x = 16'h6cba; 14'h  34: x = 16'h6c8b; 14'h  35: x = 16'h6c5d; 14'h  36: x = 16'h6c2f; 14'h  37: x = 16'h6c03; 14'h  38: x = 16'h6bd7; 14'h  39: x = 16'h6bac; 14'h  3a: x = 16'h6b82; 14'h  3b: x = 16'h6b58; 14'h  3c: x = 16'h6b2f; 14'h  3d: x = 16'h6b06; 14'h  3e: x = 16'h6adf; 14'h  3f: x = 16'h6ab7; 14'h  40: x = 16'h6a91; 14'h  41: x = 16'h6a6a; 14'h  42: x = 16'h6a45; 14'h  43: x = 16'h6a20; 14'h  44: x = 16'h69fb; 14'h  45: x = 16'h69d7; 14'h  46: x = 16'h69b3; 14'h  47: x = 16'h6990; 14'h  48: x = 16'h696d; 14'h  49: x = 16'h694b; 14'h  4a: x = 16'h6929; 14'h  4b: x = 16'h6908; 14'h  4c: x = 16'h68e7; 14'h  4d: x = 16'h68c6; 14'h  4e: x = 16'h68a6; 14'h  4f: x = 16'h6886; 14'h  50: x = 16'h6866; 14'h  51: x = 16'h6847; 14'h  52: x = 16'h6828; 14'h  53: x = 16'h680a; 14'h  54: x = 16'h67eb; 14'h  55: x = 16'h67cd; 14'h  56: x = 16'h67b0; 14'h  57: x = 16'h6793; 14'h  58: x = 16'h6776; 14'h  59: x = 16'h6759; 14'h  5a: x = 16'h673d; 14'h  5b: x = 16'h6721; 14'h  5c: x = 16'h6705; 14'h  5d: x = 16'h66e9; 14'h  5e: x = 16'h66ce; 14'h  5f: x = 16'h66b3; 14'h  60: x = 16'h6698; 14'h  61: x = 16'h667e; 14'h  62: x = 16'h6664; 14'h  63: x = 16'h664a; 14'h  64: x = 16'h6630; 14'h  65: x = 16'h6616; 14'h  66: x = 16'h65fd; 14'h  67: x = 16'h65e4; 14'h  68: x = 16'h65cb; 14'h  69: x = 16'h65b2; 14'h  6a: x = 16'h659a; 14'h  6b: x = 16'h6582; 14'h  6c: x = 16'h656a; 14'h  6d: x = 16'h6552; 14'h  6e: x = 16'h653a; 14'h  6f: x = 16'h6523; 14'h  70: x = 16'h650b; 14'h  71: x = 16'h64f4; 14'h  72: x = 16'h64dd; 14'h  73: x = 16'h64c7; 14'h  74: x = 16'h64b0; 14'h  75: x = 16'h649a; 14'h  76: x = 16'h6484; 14'h  77: x = 16'h646e; 14'h  78: x = 16'h6458; 14'h  79: x = 16'h6442; 14'h  7a: x = 16'h642d; 14'h  7b: x = 16'h6417; 14'h  7c: x = 16'h6402; 14'h  7d: x = 16'h63ed; 14'h  7e: x = 16'h63d8; 14'h  7f: x = 16'h63c3; 14'h  80: x = 16'h63af; 14'h  81: x = 16'h639a; 14'h  82: x = 16'h6386; 14'h  83: x = 16'h6372; 14'h  84: x = 16'h635e; 14'h  85: x = 16'h634a; 14'h  86: x = 16'h6336; 14'h  87: x = 16'h6322; 14'h  88: x = 16'h630f; 14'h  89: x = 16'h62fb; 14'h  8a: x = 16'h62e8; 14'h  8b: x = 16'h62d5; 14'h  8c: x = 16'h62c2; 14'h  8d: x = 16'h62af; 14'h  8e: x = 16'h629c; 14'h  8f: x = 16'h628a; 14'h  90: x = 16'h6277; 14'h  91: x = 16'h6265; 14'h  92: x = 16'h6252; 14'h  93: x = 16'h6240; 14'h  94: x = 16'h622e; 14'h  95: x = 16'h621c; 14'h  96: x = 16'h620a; 14'h  97: x = 16'h61f8; 14'h  98: x = 16'h61e7; 14'h  99: x = 16'h61d5; 14'h  9a: x = 16'h61c4; 14'h  9b: x = 16'h61b2; 14'h  9c: x = 16'h61a1; 14'h  9d: x = 16'h6190; 14'h  9e: x = 16'h617f; 14'h  9f: x = 16'h616e; 14'h  a0: x = 16'h615d; 14'h  a1: x = 16'h614c; 14'h  a2: x = 16'h613b; 14'h  a3: x = 16'h612b; 14'h  a4: x = 16'h611a; 14'h  a5: x = 16'h610a; 14'h  a6: x = 16'h60fa; 14'h  a7: x = 16'h60e9; 14'h  a8: x = 16'h60d9; 14'h  a9: x = 16'h60c9; 14'h  aa: x = 16'h60b9; 14'h  ab: x = 16'h60a9; 14'h  ac: x = 16'h6099; 14'h  ad: x = 16'h608a; 14'h  ae: x = 16'h607a; 14'h  af: x = 16'h606b; 14'h  b0: x = 16'h605b; 14'h  b1: x = 16'h604c; 14'h  b2: x = 16'h603c; 14'h  b3: x = 16'h602d; 14'h  b4: x = 16'h601e; 14'h  b5: x = 16'h600f; 14'h  b6: x = 16'h6000; 14'h  b7: x = 16'h5ff1; 14'h  b8: x = 16'h5fe2; 14'h  b9: x = 16'h5fd3; 14'h  ba: x = 16'h5fc4; 14'h  bb: x = 16'h5fb6; 14'h  bc: x = 16'h5fa7; 14'h  bd: x = 16'h5f98; 14'h  be: x = 16'h5f8a; 14'h  bf: x = 16'h5f7b; 14'h  c0: x = 16'h5f6d; 14'h  c1: x = 16'h5f5f; 14'h  c2: x = 16'h5f51; 14'h  c3: x = 16'h5f43; 14'h  c4: x = 16'h5f34; 14'h  c5: x = 16'h5f26; 14'h  c6: x = 16'h5f18; 14'h  c7: x = 16'h5f0b; 14'h  c8: x = 16'h5efd; 14'h  c9: x = 16'h5eef; 14'h  ca: x = 16'h5ee1; 14'h  cb: x = 16'h5ed4; 14'h  cc: x = 16'h5ec6; 14'h  cd: x = 16'h5eb9; 14'h  ce: x = 16'h5eab; 14'h  cf: x = 16'h5e9e; 14'h  d0: x = 16'h5e90; 14'h  d1: x = 16'h5e83; 14'h  d2: x = 16'h5e76; 14'h  d3: x = 16'h5e69; 14'h  d4: x = 16'h5e5b; 14'h  d5: x = 16'h5e4e; 14'h  d6: x = 16'h5e41; 14'h  d7: x = 16'h5e34; 14'h  d8: x = 16'h5e27; 14'h  d9: x = 16'h5e1b; 14'h  da: x = 16'h5e0e; 14'h  db: x = 16'h5e01; 14'h  dc: x = 16'h5df4; 14'h  dd: x = 16'h5de8; 14'h  de: x = 16'h5ddb; 14'h  df: x = 16'h5dce; 14'h  e0: x = 16'h5dc2; 14'h  e1: x = 16'h5db6; 14'h  e2: x = 16'h5da9; 14'h  e3: x = 16'h5d9d; 14'h  e4: x = 16'h5d90; 14'h  e5: x = 16'h5d84; 14'h  e6: x = 16'h5d78; 14'h  e7: x = 16'h5d6c; 14'h  e8: x = 16'h5d60; 14'h  e9: x = 16'h5d54; 14'h  ea: x = 16'h5d48; 14'h  eb: x = 16'h5d3c; 14'h  ec: x = 16'h5d30; 14'h  ed: x = 16'h5d24; 14'h  ee: x = 16'h5d18; 14'h  ef: x = 16'h5d0c; 14'h  f0: x = 16'h5d00; 14'h  f1: x = 16'h5cf5; 14'h  f2: x = 16'h5ce9; 14'h  f3: x = 16'h5cdd; 14'h  f4: x = 16'h5cd2; 14'h  f5: x = 16'h5cc6; 14'h  f6: x = 16'h5cbb; 14'h  f7: x = 16'h5caf; 14'h  f8: x = 16'h5ca4; 14'h  f9: x = 16'h5c98; 14'h  fa: x = 16'h5c8d; 14'h  fb: x = 16'h5c82; 14'h  fc: x = 16'h5c76; 14'h  fd: x = 16'h5c6b; 14'h  fe: x = 16'h5c60; 14'h  ff: x = 16'h5c55; 14'h 100: x = 16'h5c4a; 14'h 101: x = 16'h5c3f; 14'h 102: x = 16'h5c34; 14'h 103: x = 16'h5c29; 14'h 104: x = 16'h5c1e; 14'h 105: x = 16'h5c13; 14'h 106: x = 16'h5c08; 14'h 107: x = 16'h5bfd; 14'h 108: x = 16'h5bf2; 14'h 109: x = 16'h5be7; 14'h 10a: x = 16'h5bdd; 14'h 10b: x = 16'h5bd2; 14'h 10c: x = 16'h5bc7; 14'h 10d: x = 16'h5bbd; 14'h 10e: x = 16'h5bb2; 14'h 10f: x = 16'h5ba7; 14'h 110: x = 16'h5b9d; 14'h 111: x = 16'h5b92; 14'h 112: x = 16'h5b88; 14'h 113: x = 16'h5b7d; 14'h 114: x = 16'h5b73; 14'h 115: x = 16'h5b69; 14'h 116: x = 16'h5b5e; 14'h 117: x = 16'h5b54; 14'h 118: x = 16'h5b4a; 14'h 119: x = 16'h5b40; 14'h 11a: x = 16'h5b35; 14'h 11b: x = 16'h5b2b; 14'h 11c: x = 16'h5b21; 14'h 11d: x = 16'h5b17; 14'h 11e: x = 16'h5b0d; 14'h 11f: x = 16'h5b03; 14'h 120: x = 16'h5af9; 14'h 121: x = 16'h5aef; 14'h 122: x = 16'h5ae5; 14'h 123: x = 16'h5adb; 14'h 124: x = 16'h5ad1; 14'h 125: x = 16'h5ac7; 14'h 126: x = 16'h5abd; 14'h 127: x = 16'h5ab3; 14'h 128: x = 16'h5aaa; 14'h 129: x = 16'h5aa0; 14'h 12a: x = 16'h5a96; 14'h 12b: x = 16'h5a8c; 14'h 12c: x = 16'h5a83; 14'h 12d: x = 16'h5a79; 14'h 12e: x = 16'h5a70; 14'h 12f: x = 16'h5a66; 14'h 130: x = 16'h5a5c; 14'h 131: x = 16'h5a53; 14'h 132: x = 16'h5a49; 14'h 133: x = 16'h5a40; 14'h 134: x = 16'h5a36; 14'h 135: x = 16'h5a2d; 14'h 136: x = 16'h5a24; 14'h 137: x = 16'h5a1a; 14'h 138: x = 16'h5a11; 14'h 139: x = 16'h5a08; 14'h 13a: x = 16'h59fe; 14'h 13b: x = 16'h59f5; 14'h 13c: x = 16'h59ec; 14'h 13d: x = 16'h59e3; 14'h 13e: x = 16'h59d9; 14'h 13f: x = 16'h59d0; 14'h 140: x = 16'h59c7; 14'h 141: x = 16'h59be; 14'h 142: x = 16'h59b5; 14'h 143: x = 16'h59ac; 14'h 144: x = 16'h59a3; 14'h 145: x = 16'h599a; 14'h 146: x = 16'h5991; 14'h 147: x = 16'h5988; 14'h 148: x = 16'h597f; 14'h 149: x = 16'h5976; 14'h 14a: x = 16'h596d; 14'h 14b: x = 16'h5964; 14'h 14c: x = 16'h595b; 14'h 14d: x = 16'h5953; 14'h 14e: x = 16'h594a; 14'h 14f: x = 16'h5941; 14'h 150: x = 16'h5938; 14'h 151: x = 16'h592f; 14'h 152: x = 16'h5927; 14'h 153: x = 16'h591e; 14'h 154: x = 16'h5915; 14'h 155: x = 16'h590d; 14'h 156: x = 16'h5904; 14'h 157: x = 16'h58fc; 14'h 158: x = 16'h58f3; 14'h 159: x = 16'h58ea; 14'h 15a: x = 16'h58e2; 14'h 15b: x = 16'h58d9; 14'h 15c: x = 16'h58d1; 14'h 15d: x = 16'h58c8; 14'h 15e: x = 16'h58c0; 14'h 15f: x = 16'h58b8; 14'h 160: x = 16'h58af; 14'h 161: x = 16'h58a7; 14'h 162: x = 16'h589e; 14'h 163: x = 16'h5896; 14'h 164: x = 16'h588e; 14'h 165: x = 16'h5885; 14'h 166: x = 16'h587d; 14'h 167: x = 16'h5875; 14'h 168: x = 16'h586d; 14'h 169: x = 16'h5864; 14'h 16a: x = 16'h585c; 14'h 16b: x = 16'h5854; 14'h 16c: x = 16'h584c; 14'h 16d: x = 16'h5844; 14'h 16e: x = 16'h583c; 14'h 16f: x = 16'h5833; 14'h 170: x = 16'h582b; 14'h 171: x = 16'h5823; 14'h 172: x = 16'h581b; 14'h 173: x = 16'h5813; 14'h 174: x = 16'h580b; 14'h 175: x = 16'h5803; 14'h 176: x = 16'h57fb; 14'h 177: x = 16'h57f3; 14'h 178: x = 16'h57eb; 14'h 179: x = 16'h57e3; 14'h 17a: x = 16'h57db; 14'h 17b: x = 16'h57d4; 14'h 17c: x = 16'h57cc; 14'h 17d: x = 16'h57c4; 14'h 17e: x = 16'h57bc; 14'h 17f: x = 16'h57b4; 14'h 180: x = 16'h57ac; 14'h 181: x = 16'h57a5; 14'h 182: x = 16'h579d; 14'h 183: x = 16'h5795; 14'h 184: x = 16'h578d; 14'h 185: x = 16'h5786; 14'h 186: x = 16'h577e; 14'h 187: x = 16'h5776; 14'h 188: x = 16'h576f; 14'h 189: x = 16'h5767; 14'h 18a: x = 16'h575f; 14'h 18b: x = 16'h5758; 14'h 18c: x = 16'h5750; 14'h 18d: x = 16'h5749; 14'h 18e: x = 16'h5741; 14'h 18f: x = 16'h573a; 14'h 190: x = 16'h5732; 14'h 191: x = 16'h572b; 14'h 192: x = 16'h5723; 14'h 193: x = 16'h571c; 14'h 194: x = 16'h5714; 14'h 195: x = 16'h570d; 14'h 196: x = 16'h5705; 14'h 197: x = 16'h56fe; 14'h 198: x = 16'h56f6; 14'h 199: x = 16'h56ef; 14'h 19a: x = 16'h56e8; 14'h 19b: x = 16'h56e0; 14'h 19c: x = 16'h56d9; 14'h 19d: x = 16'h56d2; 14'h 19e: x = 16'h56ca; 14'h 19f: x = 16'h56c3; 14'h 1a0: x = 16'h56bc; 14'h 1a1: x = 16'h56b5; 14'h 1a2: x = 16'h56ad; 14'h 1a3: x = 16'h56a6; 14'h 1a4: x = 16'h569f; 14'h 1a5: x = 16'h5698; 14'h 1a6: x = 16'h5691; 14'h 1a7: x = 16'h5689; 14'h 1a8: x = 16'h5682; 14'h 1a9: x = 16'h567b; 14'h 1aa: x = 16'h5674; 14'h 1ab: x = 16'h566d; 14'h 1ac: x = 16'h5666; 14'h 1ad: x = 16'h565f; 14'h 1ae: x = 16'h5658; 14'h 1af: x = 16'h5651; 14'h 1b0: x = 16'h5649; 14'h 1b1: x = 16'h5642; 14'h 1b2: x = 16'h563b; 14'h 1b3: x = 16'h5634; 14'h 1b4: x = 16'h562d; 14'h 1b5: x = 16'h5626; 14'h 1b6: x = 16'h5620; 14'h 1b7: x = 16'h5619; 14'h 1b8: x = 16'h5612; 14'h 1b9: x = 16'h560b; 14'h 1ba: x = 16'h5604; 14'h 1bb: x = 16'h55fd; 14'h 1bc: x = 16'h55f6; 14'h 1bd: x = 16'h55ef; 14'h 1be: x = 16'h55e8; 14'h 1bf: x = 16'h55e2; 14'h 1c0: x = 16'h55db; 14'h 1c1: x = 16'h55d4; 14'h 1c2: x = 16'h55cd; 14'h 1c3: x = 16'h55c6; 14'h 1c4: x = 16'h55c0; 14'h 1c5: x = 16'h55b9; 14'h 1c6: x = 16'h55b2; 14'h 1c7: x = 16'h55ab; 14'h 1c8: x = 16'h55a5; 14'h 1c9: x = 16'h559e; 14'h 1ca: x = 16'h5597; 14'h 1cb: x = 16'h5591; 14'h 1cc: x = 16'h558a; 14'h 1cd: x = 16'h5583; 14'h 1ce: x = 16'h557d; 14'h 1cf: x = 16'h5576; 14'h 1d0: x = 16'h556f; 14'h 1d1: x = 16'h5569; 14'h 1d2: x = 16'h5562; 14'h 1d3: x = 16'h555c; 14'h 1d4: x = 16'h5555; 14'h 1d5: x = 16'h554e; 14'h 1d6: x = 16'h5548; 14'h 1d7: x = 16'h5541; 14'h 1d8: x = 16'h553b; 14'h 1d9: x = 16'h5534; 14'h 1da: x = 16'h552e; 14'h 1db: x = 16'h5527; 14'h 1dc: x = 16'h5521; 14'h 1dd: x = 16'h551a; 14'h 1de: x = 16'h5514; 14'h 1df: x = 16'h550d; 14'h 1e0: x = 16'h5507; 14'h 1e1: x = 16'h5501; 14'h 1e2: x = 16'h54fa; 14'h 1e3: x = 16'h54f4; 14'h 1e4: x = 16'h54ed; 14'h 1e5: x = 16'h54e7; 14'h 1e6: x = 16'h54e1; 14'h 1e7: x = 16'h54da; 14'h 1e8: x = 16'h54d4; 14'h 1e9: x = 16'h54ce; 14'h 1ea: x = 16'h54c7; 14'h 1eb: x = 16'h54c1; 14'h 1ec: x = 16'h54bb; 14'h 1ed: x = 16'h54b4; 14'h 1ee: x = 16'h54ae; 14'h 1ef: x = 16'h54a8; 14'h 1f0: x = 16'h54a2; 14'h 1f1: x = 16'h549b; 14'h 1f2: x = 16'h5495; 14'h 1f3: x = 16'h548f; 14'h 1f4: x = 16'h5489; 14'h 1f5: x = 16'h5483; 14'h 1f6: x = 16'h547c; 14'h 1f7: x = 16'h5476; 14'h 1f8: x = 16'h5470; 14'h 1f9: x = 16'h546a; 14'h 1fa: x = 16'h5464; 14'h 1fb: x = 16'h545e; 14'h 1fc: x = 16'h5458; 14'h 1fd: x = 16'h5451; 14'h 1fe: x = 16'h544b; 14'h 1ff: x = 16'h5445; 14'h 200: x = 16'h543f; 14'h 201: x = 16'h5439; 14'h 202: x = 16'h5433; 14'h 203: x = 16'h542d; 14'h 204: x = 16'h5427; 14'h 205: x = 16'h5421; 14'h 206: x = 16'h541b; 14'h 207: x = 16'h5415; 14'h 208: x = 16'h540f; 14'h 209: x = 16'h5409; 14'h 20a: x = 16'h5403; 14'h 20b: x = 16'h53fd; 14'h 20c: x = 16'h53f7; 14'h 20d: x = 16'h53f1; 14'h 20e: x = 16'h53eb; 14'h 20f: x = 16'h53e5; 14'h 210: x = 16'h53df; 14'h 211: x = 16'h53d9; 14'h 212: x = 16'h53d3; 14'h 213: x = 16'h53cd; 14'h 214: x = 16'h53c8; 14'h 215: x = 16'h53c2; 14'h 216: x = 16'h53bc; 14'h 217: x = 16'h53b6; 14'h 218: x = 16'h53b0; 14'h 219: x = 16'h53aa; 14'h 21a: x = 16'h53a4; 14'h 21b: x = 16'h539f; 14'h 21c: x = 16'h5399; 14'h 21d: x = 16'h5393; 14'h 21e: x = 16'h538d; 14'h 21f: x = 16'h5387; 14'h 220: x = 16'h5382; 14'h 221: x = 16'h537c; 14'h 222: x = 16'h5376; 14'h 223: x = 16'h5370; 14'h 224: x = 16'h536b; 14'h 225: x = 16'h5365; 14'h 226: x = 16'h535f; 14'h 227: x = 16'h535a; 14'h 228: x = 16'h5354; 14'h 229: x = 16'h534e; 14'h 22a: x = 16'h5348; 14'h 22b: x = 16'h5343; 14'h 22c: x = 16'h533d; 14'h 22d: x = 16'h5337; 14'h 22e: x = 16'h5332; 14'h 22f: x = 16'h532c; 14'h 230: x = 16'h5326; 14'h 231: x = 16'h5321; 14'h 232: x = 16'h531b; 14'h 233: x = 16'h5316; 14'h 234: x = 16'h5310; 14'h 235: x = 16'h530a; 14'h 236: x = 16'h5305; 14'h 237: x = 16'h52ff; 14'h 238: x = 16'h52fa; 14'h 239: x = 16'h52f4; 14'h 23a: x = 16'h52ef; 14'h 23b: x = 16'h52e9; 14'h 23c: x = 16'h52e4; 14'h 23d: x = 16'h52de; 14'h 23e: x = 16'h52d8; 14'h 23f: x = 16'h52d3; 14'h 240: x = 16'h52cd; 14'h 241: x = 16'h52c8; 14'h 242: x = 16'h52c3; 14'h 243: x = 16'h52bd; 14'h 244: x = 16'h52b8; 14'h 245: x = 16'h52b2; 14'h 246: x = 16'h52ad; 14'h 247: x = 16'h52a7; 14'h 248: x = 16'h52a2; 14'h 249: x = 16'h529c; 14'h 24a: x = 16'h5297; 14'h 24b: x = 16'h5292; 14'h 24c: x = 16'h528c; 14'h 24d: x = 16'h5287; 14'h 24e: x = 16'h5281; 14'h 24f: x = 16'h527c; 14'h 250: x = 16'h5277; 14'h 251: x = 16'h5271; 14'h 252: x = 16'h526c; 14'h 253: x = 16'h5266; 14'h 254: x = 16'h5261; 14'h 255: x = 16'h525c; 14'h 256: x = 16'h5256; 14'h 257: x = 16'h5251; 14'h 258: x = 16'h524c; 14'h 259: x = 16'h5247; 14'h 25a: x = 16'h5241; 14'h 25b: x = 16'h523c; 14'h 25c: x = 16'h5237; 14'h 25d: x = 16'h5231; 14'h 25e: x = 16'h522c; 14'h 25f: x = 16'h5227; 14'h 260: x = 16'h5222; 14'h 261: x = 16'h521c; 14'h 262: x = 16'h5217; 14'h 263: x = 16'h5212; 14'h 264: x = 16'h520d; 14'h 265: x = 16'h5207; 14'h 266: x = 16'h5202; 14'h 267: x = 16'h51fd; 14'h 268: x = 16'h51f8; 14'h 269: x = 16'h51f3; 14'h 26a: x = 16'h51ed; 14'h 26b: x = 16'h51e8; 14'h 26c: x = 16'h51e3; 14'h 26d: x = 16'h51de; 14'h 26e: x = 16'h51d9; 14'h 26f: x = 16'h51d4; 14'h 270: x = 16'h51cf; 14'h 271: x = 16'h51c9; 14'h 272: x = 16'h51c4; 14'h 273: x = 16'h51bf; 14'h 274: x = 16'h51ba; 14'h 275: x = 16'h51b5; 14'h 276: x = 16'h51b0; 14'h 277: x = 16'h51ab; 14'h 278: x = 16'h51a6; 14'h 279: x = 16'h51a1; 14'h 27a: x = 16'h519c; 14'h 27b: x = 16'h5196; 14'h 27c: x = 16'h5191; 14'h 27d: x = 16'h518c; 14'h 27e: x = 16'h5187; 14'h 27f: x = 16'h5182; 14'h 280: x = 16'h517d; 14'h 281: x = 16'h5178; 14'h 282: x = 16'h5173; 14'h 283: x = 16'h516e; 14'h 284: x = 16'h5169; 14'h 285: x = 16'h5164; 14'h 286: x = 16'h515f; 14'h 287: x = 16'h515a; 14'h 288: x = 16'h5155; 14'h 289: x = 16'h5150; 14'h 28a: x = 16'h514b; 14'h 28b: x = 16'h5146; 14'h 28c: x = 16'h5141; 14'h 28d: x = 16'h513c; 14'h 28e: x = 16'h5138; 14'h 28f: x = 16'h5133; 14'h 290: x = 16'h512e; 14'h 291: x = 16'h5129; 14'h 292: x = 16'h5124; 14'h 293: x = 16'h511f; 14'h 294: x = 16'h511a; 14'h 295: x = 16'h5115; 14'h 296: x = 16'h5110; 14'h 297: x = 16'h510b; 14'h 298: x = 16'h5107; 14'h 299: x = 16'h5102; 14'h 29a: x = 16'h50fd; 14'h 29b: x = 16'h50f8; 14'h 29c: x = 16'h50f3; 14'h 29d: x = 16'h50ee; 14'h 29e: x = 16'h50e9; 14'h 29f: x = 16'h50e5; 14'h 2a0: x = 16'h50e0; 14'h 2a1: x = 16'h50db; 14'h 2a2: x = 16'h50d6; 14'h 2a3: x = 16'h50d1; 14'h 2a4: x = 16'h50cc; 14'h 2a5: x = 16'h50c8; 14'h 2a6: x = 16'h50c3; 14'h 2a7: x = 16'h50be; 14'h 2a8: x = 16'h50b9; 14'h 2a9: x = 16'h50b5; 14'h 2aa: x = 16'h50b0; 14'h 2ab: x = 16'h50ab; 14'h 2ac: x = 16'h50a6; 14'h 2ad: x = 16'h50a2; 14'h 2ae: x = 16'h509d; 14'h 2af: x = 16'h5098; 14'h 2b0: x = 16'h5093; 14'h 2b1: x = 16'h508f; 14'h 2b2: x = 16'h508a; 14'h 2b3: x = 16'h5085; 14'h 2b4: x = 16'h5080; 14'h 2b5: x = 16'h507c; 14'h 2b6: x = 16'h5077; 14'h 2b7: x = 16'h5072; 14'h 2b8: x = 16'h506e; 14'h 2b9: x = 16'h5069; 14'h 2ba: x = 16'h5064; 14'h 2bb: x = 16'h5060; 14'h 2bc: x = 16'h505b; 14'h 2bd: x = 16'h5056; 14'h 2be: x = 16'h5052; 14'h 2bf: x = 16'h504d; 14'h 2c0: x = 16'h5048; 14'h 2c1: x = 16'h5044; 14'h 2c2: x = 16'h503f; 14'h 2c3: x = 16'h503a; 14'h 2c4: x = 16'h5036; 14'h 2c5: x = 16'h5031; 14'h 2c6: x = 16'h502d; 14'h 2c7: x = 16'h5028; 14'h 2c8: x = 16'h5023; 14'h 2c9: x = 16'h501f; 14'h 2ca: x = 16'h501a; 14'h 2cb: x = 16'h5016; 14'h 2cc: x = 16'h5011; 14'h 2cd: x = 16'h500d; 14'h 2ce: x = 16'h5008; 14'h 2cf: x = 16'h5003; 14'h 2d0: x = 16'h4fff; 14'h 2d1: x = 16'h4ffa; 14'h 2d2: x = 16'h4ff6; 14'h 2d3: x = 16'h4ff1; 14'h 2d4: x = 16'h4fed; 14'h 2d5: x = 16'h4fe8; 14'h 2d6: x = 16'h4fe4; 14'h 2d7: x = 16'h4fdf; 14'h 2d8: x = 16'h4fdb; 14'h 2d9: x = 16'h4fd6; 14'h 2da: x = 16'h4fd2; 14'h 2db: x = 16'h4fcd; 14'h 2dc: x = 16'h4fc9; 14'h 2dd: x = 16'h4fc4; 14'h 2de: x = 16'h4fc0; 14'h 2df: x = 16'h4fbb; 14'h 2e0: x = 16'h4fb7; 14'h 2e1: x = 16'h4fb2; 14'h 2e2: x = 16'h4fae; 14'h 2e3: x = 16'h4fa9; 14'h 2e4: x = 16'h4fa5; 14'h 2e5: x = 16'h4fa0; 14'h 2e6: x = 16'h4f9c; 14'h 2e7: x = 16'h4f98; 14'h 2e8: x = 16'h4f93; 14'h 2e9: x = 16'h4f8f; 14'h 2ea: x = 16'h4f8a; 14'h 2eb: x = 16'h4f86; 14'h 2ec: x = 16'h4f81; 14'h 2ed: x = 16'h4f7d; 14'h 2ee: x = 16'h4f79; 14'h 2ef: x = 16'h4f74; 14'h 2f0: x = 16'h4f70; 14'h 2f1: x = 16'h4f6b; 14'h 2f2: x = 16'h4f67; 14'h 2f3: x = 16'h4f63; 14'h 2f4: x = 16'h4f5e; 14'h 2f5: x = 16'h4f5a; 14'h 2f6: x = 16'h4f56; 14'h 2f7: x = 16'h4f51; 14'h 2f8: x = 16'h4f4d; 14'h 2f9: x = 16'h4f49; 14'h 2fa: x = 16'h4f44; 14'h 2fb: x = 16'h4f40; 14'h 2fc: x = 16'h4f3c; 14'h 2fd: x = 16'h4f37; 14'h 2fe: x = 16'h4f33; 14'h 2ff: x = 16'h4f2f; 14'h 300: x = 16'h4f2a; 14'h 301: x = 16'h4f26; 14'h 302: x = 16'h4f22; 14'h 303: x = 16'h4f1d; 14'h 304: x = 16'h4f19; 14'h 305: x = 16'h4f15; 14'h 306: x = 16'h4f11; 14'h 307: x = 16'h4f0c; 14'h 308: x = 16'h4f08; 14'h 309: x = 16'h4f04; 14'h 30a: x = 16'h4eff; 14'h 30b: x = 16'h4efb; 14'h 30c: x = 16'h4ef7; 14'h 30d: x = 16'h4ef3; 14'h 30e: x = 16'h4eee; 14'h 30f: x = 16'h4eea; 14'h 310: x = 16'h4ee6; 14'h 311: x = 16'h4ee2; 14'h 312: x = 16'h4edd; 14'h 313: x = 16'h4ed9; 14'h 314: x = 16'h4ed5; 14'h 315: x = 16'h4ed1; 14'h 316: x = 16'h4ecd; 14'h 317: x = 16'h4ec8; 14'h 318: x = 16'h4ec4; 14'h 319: x = 16'h4ec0; 14'h 31a: x = 16'h4ebc; 14'h 31b: x = 16'h4eb8; 14'h 31c: x = 16'h4eb3; 14'h 31d: x = 16'h4eaf; 14'h 31e: x = 16'h4eab; 14'h 31f: x = 16'h4ea7; 14'h 320: x = 16'h4ea3; 14'h 321: x = 16'h4e9e; 14'h 322: x = 16'h4e9a; 14'h 323: x = 16'h4e96; 14'h 324: x = 16'h4e92; 14'h 325: x = 16'h4e8e; 14'h 326: x = 16'h4e8a; 14'h 327: x = 16'h4e86; 14'h 328: x = 16'h4e81; 14'h 329: x = 16'h4e7d; 14'h 32a: x = 16'h4e79; 14'h 32b: x = 16'h4e75; 14'h 32c: x = 16'h4e71; 14'h 32d: x = 16'h4e6d; 14'h 32e: x = 16'h4e69; 14'h 32f: x = 16'h4e65; 14'h 330: x = 16'h4e61; 14'h 331: x = 16'h4e5c; 14'h 332: x = 16'h4e58; 14'h 333: x = 16'h4e54; 14'h 334: x = 16'h4e50; 14'h 335: x = 16'h4e4c; 14'h 336: x = 16'h4e48; 14'h 337: x = 16'h4e44; 14'h 338: x = 16'h4e40; 14'h 339: x = 16'h4e3c; 14'h 33a: x = 16'h4e38; 14'h 33b: x = 16'h4e34; 14'h 33c: x = 16'h4e30; 14'h 33d: x = 16'h4e2c; 14'h 33e: x = 16'h4e28; 14'h 33f: x = 16'h4e24; 14'h 340: x = 16'h4e1f; 14'h 341: x = 16'h4e1b; 14'h 342: x = 16'h4e17; 14'h 343: x = 16'h4e13; 14'h 344: x = 16'h4e0f; 14'h 345: x = 16'h4e0b; 14'h 346: x = 16'h4e07; 14'h 347: x = 16'h4e03; 14'h 348: x = 16'h4dff; 14'h 349: x = 16'h4dfb; 14'h 34a: x = 16'h4df7; 14'h 34b: x = 16'h4df3; 14'h 34c: x = 16'h4def; 14'h 34d: x = 16'h4deb; 14'h 34e: x = 16'h4de7; 14'h 34f: x = 16'h4de3; 14'h 350: x = 16'h4ddf; 14'h 351: x = 16'h4ddc; 14'h 352: x = 16'h4dd8; 14'h 353: x = 16'h4dd4; 14'h 354: x = 16'h4dd0; 14'h 355: x = 16'h4dcc; 14'h 356: x = 16'h4dc8; 14'h 357: x = 16'h4dc4; 14'h 358: x = 16'h4dc0; 14'h 359: x = 16'h4dbc; 14'h 35a: x = 16'h4db8; 14'h 35b: x = 16'h4db4; 14'h 35c: x = 16'h4db0; 14'h 35d: x = 16'h4dac; 14'h 35e: x = 16'h4da8; 14'h 35f: x = 16'h4da4; 14'h 360: x = 16'h4da0; 14'h 361: x = 16'h4d9d; 14'h 362: x = 16'h4d99; 14'h 363: x = 16'h4d95; 14'h 364: x = 16'h4d91; 14'h 365: x = 16'h4d8d; 14'h 366: x = 16'h4d89; 14'h 367: x = 16'h4d85; 14'h 368: x = 16'h4d81; 14'h 369: x = 16'h4d7d; 14'h 36a: x = 16'h4d7a; 14'h 36b: x = 16'h4d76; 14'h 36c: x = 16'h4d72; 14'h 36d: x = 16'h4d6e; 14'h 36e: x = 16'h4d6a; 14'h 36f: x = 16'h4d66; 14'h 370: x = 16'h4d62; 14'h 371: x = 16'h4d5f; 14'h 372: x = 16'h4d5b; 14'h 373: x = 16'h4d57; 14'h 374: x = 16'h4d53; 14'h 375: x = 16'h4d4f; 14'h 376: x = 16'h4d4b; 14'h 377: x = 16'h4d48; 14'h 378: x = 16'h4d44; 14'h 379: x = 16'h4d40; 14'h 37a: x = 16'h4d3c; 14'h 37b: x = 16'h4d38; 14'h 37c: x = 16'h4d34; 14'h 37d: x = 16'h4d31; 14'h 37e: x = 16'h4d2d; 14'h 37f: x = 16'h4d29; 14'h 380: x = 16'h4d25; 14'h 381: x = 16'h4d21; 14'h 382: x = 16'h4d1e; 14'h 383: x = 16'h4d1a; 14'h 384: x = 16'h4d16; 14'h 385: x = 16'h4d12; 14'h 386: x = 16'h4d0f; 14'h 387: x = 16'h4d0b; 14'h 388: x = 16'h4d07; 14'h 389: x = 16'h4d03; 14'h 38a: x = 16'h4d00; 14'h 38b: x = 16'h4cfc; 14'h 38c: x = 16'h4cf8; 14'h 38d: x = 16'h4cf4; 14'h 38e: x = 16'h4cf1; 14'h 38f: x = 16'h4ced; 14'h 390: x = 16'h4ce9; 14'h 391: x = 16'h4ce5; 14'h 392: x = 16'h4ce2; 14'h 393: x = 16'h4cde; 14'h 394: x = 16'h4cda; 14'h 395: x = 16'h4cd6; 14'h 396: x = 16'h4cd3; 14'h 397: x = 16'h4ccf; 14'h 398: x = 16'h4ccb; 14'h 399: x = 16'h4cc8; 14'h 39a: x = 16'h4cc4; 14'h 39b: x = 16'h4cc0; 14'h 39c: x = 16'h4cbc; 14'h 39d: x = 16'h4cb9; 14'h 39e: x = 16'h4cb5; 14'h 39f: x = 16'h4cb1; 14'h 3a0: x = 16'h4cae; 14'h 3a1: x = 16'h4caa; 14'h 3a2: x = 16'h4ca6; 14'h 3a3: x = 16'h4ca3; 14'h 3a4: x = 16'h4c9f; 14'h 3a5: x = 16'h4c9b; 14'h 3a6: x = 16'h4c98; 14'h 3a7: x = 16'h4c94; 14'h 3a8: x = 16'h4c90; 14'h 3a9: x = 16'h4c8d; 14'h 3aa: x = 16'h4c89; 14'h 3ab: x = 16'h4c85; 14'h 3ac: x = 16'h4c82; 14'h 3ad: x = 16'h4c7e; 14'h 3ae: x = 16'h4c7a; 14'h 3af: x = 16'h4c77; 14'h 3b0: x = 16'h4c73; 14'h 3b1: x = 16'h4c6f; 14'h 3b2: x = 16'h4c6c; 14'h 3b3: x = 16'h4c68; 14'h 3b4: x = 16'h4c65; 14'h 3b5: x = 16'h4c61; 14'h 3b6: x = 16'h4c5d; 14'h 3b7: x = 16'h4c5a; 14'h 3b8: x = 16'h4c56; 14'h 3b9: x = 16'h4c53; 14'h 3ba: x = 16'h4c4f; 14'h 3bb: x = 16'h4c4b; 14'h 3bc: x = 16'h4c48; 14'h 3bd: x = 16'h4c44; 14'h 3be: x = 16'h4c41; 14'h 3bf: x = 16'h4c3d; 14'h 3c0: x = 16'h4c39; 14'h 3c1: x = 16'h4c36; 14'h 3c2: x = 16'h4c32; 14'h 3c3: x = 16'h4c2f; 14'h 3c4: x = 16'h4c2b; 14'h 3c5: x = 16'h4c28; 14'h 3c6: x = 16'h4c24; 14'h 3c7: x = 16'h4c20; 14'h 3c8: x = 16'h4c1d; 14'h 3c9: x = 16'h4c19; 14'h 3ca: x = 16'h4c16; 14'h 3cb: x = 16'h4c12; 14'h 3cc: x = 16'h4c0f; 14'h 3cd: x = 16'h4c0b; 14'h 3ce: x = 16'h4c08; 14'h 3cf: x = 16'h4c04; 14'h 3d0: x = 16'h4c00; 14'h 3d1: x = 16'h4bfd; 14'h 3d2: x = 16'h4bf9; 14'h 3d3: x = 16'h4bf6; 14'h 3d4: x = 16'h4bf2; 14'h 3d5: x = 16'h4bef; 14'h 3d6: x = 16'h4beb; 14'h 3d7: x = 16'h4be8; 14'h 3d8: x = 16'h4be4; 14'h 3d9: x = 16'h4be1; 14'h 3da: x = 16'h4bdd; 14'h 3db: x = 16'h4bda; 14'h 3dc: x = 16'h4bd6; 14'h 3dd: x = 16'h4bd3; 14'h 3de: x = 16'h4bcf; 14'h 3df: x = 16'h4bcc; 14'h 3e0: x = 16'h4bc8; 14'h 3e1: x = 16'h4bc5; 14'h 3e2: x = 16'h4bc1; 14'h 3e3: x = 16'h4bbe; 14'h 3e4: x = 16'h4bba; 14'h 3e5: x = 16'h4bb7; 14'h 3e6: x = 16'h4bb3; 14'h 3e7: x = 16'h4bb0; 14'h 3e8: x = 16'h4bad; 14'h 3e9: x = 16'h4ba9; 14'h 3ea: x = 16'h4ba6; 14'h 3eb: x = 16'h4ba2; 14'h 3ec: x = 16'h4b9f; 14'h 3ed: x = 16'h4b9b; 14'h 3ee: x = 16'h4b98; 14'h 3ef: x = 16'h4b94; 14'h 3f0: x = 16'h4b91; 14'h 3f1: x = 16'h4b8d; 14'h 3f2: x = 16'h4b8a; 14'h 3f3: x = 16'h4b87; 14'h 3f4: x = 16'h4b83; 14'h 3f5: x = 16'h4b80; 14'h 3f6: x = 16'h4b7c; 14'h 3f7: x = 16'h4b79; 14'h 3f8: x = 16'h4b75; 14'h 3f9: x = 16'h4b72; 14'h 3fa: x = 16'h4b6f; 14'h 3fb: x = 16'h4b6b; 14'h 3fc: x = 16'h4b68; 14'h 3fd: x = 16'h4b64; 14'h 3fe: x = 16'h4b61; 14'h 3ff: x = 16'h4b5e; 14'h 400: x = 16'h4b5a; 14'h 401: x = 16'h4b57; 14'h 402: x = 16'h4b53; 14'h 403: x = 16'h4b50; 14'h 404: x = 16'h4b4d; 14'h 405: x = 16'h4b49; 14'h 406: x = 16'h4b46; 14'h 407: x = 16'h4b42; 14'h 408: x = 16'h4b3f; 14'h 409: x = 16'h4b3c; 14'h 40a: x = 16'h4b38; 14'h 40b: x = 16'h4b35; 14'h 40c: x = 16'h4b32; 14'h 40d: x = 16'h4b2e; 14'h 40e: x = 16'h4b2b; 14'h 40f: x = 16'h4b28; 14'h 410: x = 16'h4b24; 14'h 411: x = 16'h4b21; 14'h 412: x = 16'h4b1d; 14'h 413: x = 16'h4b1a; 14'h 414: x = 16'h4b17; 14'h 415: x = 16'h4b13; 14'h 416: x = 16'h4b10; 14'h 417: x = 16'h4b0d; 14'h 418: x = 16'h4b09; 14'h 419: x = 16'h4b06; 14'h 41a: x = 16'h4b03; 14'h 41b: x = 16'h4aff; 14'h 41c: x = 16'h4afc; 14'h 41d: x = 16'h4af9; 14'h 41e: x = 16'h4af5; 14'h 41f: x = 16'h4af2; 14'h 420: x = 16'h4aef; 14'h 421: x = 16'h4aec; 14'h 422: x = 16'h4ae8; 14'h 423: x = 16'h4ae5; 14'h 424: x = 16'h4ae2; 14'h 425: x = 16'h4ade; 14'h 426: x = 16'h4adb; 14'h 427: x = 16'h4ad8; 14'h 428: x = 16'h4ad4; 14'h 429: x = 16'h4ad1; 14'h 42a: x = 16'h4ace; 14'h 42b: x = 16'h4acb; 14'h 42c: x = 16'h4ac7; 14'h 42d: x = 16'h4ac4; 14'h 42e: x = 16'h4ac1; 14'h 42f: x = 16'h4abd; 14'h 430: x = 16'h4aba; 14'h 431: x = 16'h4ab7; 14'h 432: x = 16'h4ab4; 14'h 433: x = 16'h4ab0; 14'h 434: x = 16'h4aad; 14'h 435: x = 16'h4aaa; 14'h 436: x = 16'h4aa7; 14'h 437: x = 16'h4aa3; 14'h 438: x = 16'h4aa0; 14'h 439: x = 16'h4a9d; 14'h 43a: x = 16'h4a9a; 14'h 43b: x = 16'h4a96; 14'h 43c: x = 16'h4a93; 14'h 43d: x = 16'h4a90; 14'h 43e: x = 16'h4a8d; 14'h 43f: x = 16'h4a89; 14'h 440: x = 16'h4a86; 14'h 441: x = 16'h4a83; 14'h 442: x = 16'h4a80; 14'h 443: x = 16'h4a7c; 14'h 444: x = 16'h4a79; 14'h 445: x = 16'h4a76; 14'h 446: x = 16'h4a73; 14'h 447: x = 16'h4a70; 14'h 448: x = 16'h4a6c; 14'h 449: x = 16'h4a69; 14'h 44a: x = 16'h4a66; 14'h 44b: x = 16'h4a63; 14'h 44c: x = 16'h4a5f; 14'h 44d: x = 16'h4a5c; 14'h 44e: x = 16'h4a59; 14'h 44f: x = 16'h4a56; 14'h 450: x = 16'h4a53; 14'h 451: x = 16'h4a50; 14'h 452: x = 16'h4a4c; 14'h 453: x = 16'h4a49; 14'h 454: x = 16'h4a46; 14'h 455: x = 16'h4a43; 14'h 456: x = 16'h4a40; 14'h 457: x = 16'h4a3c; 14'h 458: x = 16'h4a39; 14'h 459: x = 16'h4a36; 14'h 45a: x = 16'h4a33; 14'h 45b: x = 16'h4a30; 14'h 45c: x = 16'h4a2d; 14'h 45d: x = 16'h4a29; 14'h 45e: x = 16'h4a26; 14'h 45f: x = 16'h4a23; 14'h 460: x = 16'h4a20; 14'h 461: x = 16'h4a1d; 14'h 462: x = 16'h4a1a; 14'h 463: x = 16'h4a16; 14'h 464: x = 16'h4a13; 14'h 465: x = 16'h4a10; 14'h 466: x = 16'h4a0d; 14'h 467: x = 16'h4a0a; 14'h 468: x = 16'h4a07; 14'h 469: x = 16'h4a04; 14'h 46a: x = 16'h4a00; 14'h 46b: x = 16'h49fd; 14'h 46c: x = 16'h49fa; 14'h 46d: x = 16'h49f7; 14'h 46e: x = 16'h49f4; 14'h 46f: x = 16'h49f1; 14'h 470: x = 16'h49ee; 14'h 471: x = 16'h49eb; 14'h 472: x = 16'h49e7; 14'h 473: x = 16'h49e4; 14'h 474: x = 16'h49e1; 14'h 475: x = 16'h49de; 14'h 476: x = 16'h49db; 14'h 477: x = 16'h49d8; 14'h 478: x = 16'h49d5; 14'h 479: x = 16'h49d2; 14'h 47a: x = 16'h49cf; 14'h 47b: x = 16'h49cb; 14'h 47c: x = 16'h49c8; 14'h 47d: x = 16'h49c5; 14'h 47e: x = 16'h49c2; 14'h 47f: x = 16'h49bf; 14'h 480: x = 16'h49bc; 14'h 481: x = 16'h49b9; 14'h 482: x = 16'h49b6; 14'h 483: x = 16'h49b3; 14'h 484: x = 16'h49b0; 14'h 485: x = 16'h49ad; 14'h 486: x = 16'h49aa; 14'h 487: x = 16'h49a6; 14'h 488: x = 16'h49a3; 14'h 489: x = 16'h49a0; 14'h 48a: x = 16'h499d; 14'h 48b: x = 16'h499a; 14'h 48c: x = 16'h4997; 14'h 48d: x = 16'h4994; 14'h 48e: x = 16'h4991; 14'h 48f: x = 16'h498e; 14'h 490: x = 16'h498b; 14'h 491: x = 16'h4988; 14'h 492: x = 16'h4985; 14'h 493: x = 16'h4982; 14'h 494: x = 16'h497f; 14'h 495: x = 16'h497c; 14'h 496: x = 16'h4979; 14'h 497: x = 16'h4976; 14'h 498: x = 16'h4973; 14'h 499: x = 16'h4970; 14'h 49a: x = 16'h496c; 14'h 49b: x = 16'h4969; 14'h 49c: x = 16'h4966; 14'h 49d: x = 16'h4963; 14'h 49e: x = 16'h4960; 14'h 49f: x = 16'h495d; 14'h 4a0: x = 16'h495a; 14'h 4a1: x = 16'h4957; 14'h 4a2: x = 16'h4954; 14'h 4a3: x = 16'h4951; 14'h 4a4: x = 16'h494e; 14'h 4a5: x = 16'h494b; 14'h 4a6: x = 16'h4948; 14'h 4a7: x = 16'h4945; 14'h 4a8: x = 16'h4942; 14'h 4a9: x = 16'h493f; 14'h 4aa: x = 16'h493c; 14'h 4ab: x = 16'h4939; 14'h 4ac: x = 16'h4936; 14'h 4ad: x = 16'h4933; 14'h 4ae: x = 16'h4930; 14'h 4af: x = 16'h492d; 14'h 4b0: x = 16'h492a; 14'h 4b1: x = 16'h4927; 14'h 4b2: x = 16'h4924; 14'h 4b3: x = 16'h4921; 14'h 4b4: x = 16'h491e; 14'h 4b5: x = 16'h491b; 14'h 4b6: x = 16'h4918; 14'h 4b7: x = 16'h4915; 14'h 4b8: x = 16'h4912; 14'h 4b9: x = 16'h4910; 14'h 4ba: x = 16'h490d; 14'h 4bb: x = 16'h490a; 14'h 4bc: x = 16'h4907; 14'h 4bd: x = 16'h4904; 14'h 4be: x = 16'h4901; 14'h 4bf: x = 16'h48fe; 14'h 4c0: x = 16'h48fb; 14'h 4c1: x = 16'h48f8; 14'h 4c2: x = 16'h48f5; 14'h 4c3: x = 16'h48f2; 14'h 4c4: x = 16'h48ef; 14'h 4c5: x = 16'h48ec; 14'h 4c6: x = 16'h48e9; 14'h 4c7: x = 16'h48e6; 14'h 4c8: x = 16'h48e3; 14'h 4c9: x = 16'h48e0; 14'h 4ca: x = 16'h48dd; 14'h 4cb: x = 16'h48da; 14'h 4cc: x = 16'h48d7; 14'h 4cd: x = 16'h48d5; 14'h 4ce: x = 16'h48d2; 14'h 4cf: x = 16'h48cf; 14'h 4d0: x = 16'h48cc; 14'h 4d1: x = 16'h48c9; 14'h 4d2: x = 16'h48c6; 14'h 4d3: x = 16'h48c3; 14'h 4d4: x = 16'h48c0; 14'h 4d5: x = 16'h48bd; 14'h 4d6: x = 16'h48ba; 14'h 4d7: x = 16'h48b7; 14'h 4d8: x = 16'h48b4; 14'h 4d9: x = 16'h48b2; 14'h 4da: x = 16'h48af; 14'h 4db: x = 16'h48ac; 14'h 4dc: x = 16'h48a9; 14'h 4dd: x = 16'h48a6; 14'h 4de: x = 16'h48a3; 14'h 4df: x = 16'h48a0; 14'h 4e0: x = 16'h489d; 14'h 4e1: x = 16'h489a; 14'h 4e2: x = 16'h4897; 14'h 4e3: x = 16'h4895; 14'h 4e4: x = 16'h4892; 14'h 4e5: x = 16'h488f; 14'h 4e6: x = 16'h488c; 14'h 4e7: x = 16'h4889; 14'h 4e8: x = 16'h4886; 14'h 4e9: x = 16'h4883; 14'h 4ea: x = 16'h4880; 14'h 4eb: x = 16'h487e; 14'h 4ec: x = 16'h487b; 14'h 4ed: x = 16'h4878; 14'h 4ee: x = 16'h4875; 14'h 4ef: x = 16'h4872; 14'h 4f0: x = 16'h486f; 14'h 4f1: x = 16'h486c; 14'h 4f2: x = 16'h4869; 14'h 4f3: x = 16'h4867; 14'h 4f4: x = 16'h4864; 14'h 4f5: x = 16'h4861; 14'h 4f6: x = 16'h485e; 14'h 4f7: x = 16'h485b; 14'h 4f8: x = 16'h4858; 14'h 4f9: x = 16'h4856; 14'h 4fa: x = 16'h4853; 14'h 4fb: x = 16'h4850; 14'h 4fc: x = 16'h484d; 14'h 4fd: x = 16'h484a; 14'h 4fe: x = 16'h4847; 14'h 4ff: x = 16'h4844; 14'h 500: x = 16'h4842; 14'h 501: x = 16'h483f; 14'h 502: x = 16'h483c; 14'h 503: x = 16'h4839; 14'h 504: x = 16'h4836; 14'h 505: x = 16'h4833; 14'h 506: x = 16'h4831; 14'h 507: x = 16'h482e; 14'h 508: x = 16'h482b; 14'h 509: x = 16'h4828; 14'h 50a: x = 16'h4825; 14'h 50b: x = 16'h4823; 14'h 50c: x = 16'h4820; 14'h 50d: x = 16'h481d; 14'h 50e: x = 16'h481a; 14'h 50f: x = 16'h4817; 14'h 510: x = 16'h4815; 14'h 511: x = 16'h4812; 14'h 512: x = 16'h480f; 14'h 513: x = 16'h480c; 14'h 514: x = 16'h4809; 14'h 515: x = 16'h4806; 14'h 516: x = 16'h4804; 14'h 517: x = 16'h4801; 14'h 518: x = 16'h47fe; 14'h 519: x = 16'h47fb; 14'h 51a: x = 16'h47f9; 14'h 51b: x = 16'h47f6; 14'h 51c: x = 16'h47f3; 14'h 51d: x = 16'h47f0; 14'h 51e: x = 16'h47ed; 14'h 51f: x = 16'h47eb; 14'h 520: x = 16'h47e8; 14'h 521: x = 16'h47e5; 14'h 522: x = 16'h47e2; 14'h 523: x = 16'h47e0; 14'h 524: x = 16'h47dd; 14'h 525: x = 16'h47da; 14'h 526: x = 16'h47d7; 14'h 527: x = 16'h47d4; 14'h 528: x = 16'h47d2; 14'h 529: x = 16'h47cf; 14'h 52a: x = 16'h47cc; 14'h 52b: x = 16'h47c9; 14'h 52c: x = 16'h47c7; 14'h 52d: x = 16'h47c4; 14'h 52e: x = 16'h47c1; 14'h 52f: x = 16'h47be; 14'h 530: x = 16'h47bc; 14'h 531: x = 16'h47b9; 14'h 532: x = 16'h47b6; 14'h 533: x = 16'h47b3; 14'h 534: x = 16'h47b1; 14'h 535: x = 16'h47ae; 14'h 536: x = 16'h47ab; 14'h 537: x = 16'h47a8; 14'h 538: x = 16'h47a6; 14'h 539: x = 16'h47a3; 14'h 53a: x = 16'h47a0; 14'h 53b: x = 16'h479d; 14'h 53c: x = 16'h479b; 14'h 53d: x = 16'h4798; 14'h 53e: x = 16'h4795; 14'h 53f: x = 16'h4792; 14'h 540: x = 16'h4790; 14'h 541: x = 16'h478d; 14'h 542: x = 16'h478a; 14'h 543: x = 16'h4788; 14'h 544: x = 16'h4785; 14'h 545: x = 16'h4782; 14'h 546: x = 16'h477f; 14'h 547: x = 16'h477d; 14'h 548: x = 16'h477a; 14'h 549: x = 16'h4777; 14'h 54a: x = 16'h4775; 14'h 54b: x = 16'h4772; 14'h 54c: x = 16'h476f; 14'h 54d: x = 16'h476c; 14'h 54e: x = 16'h476a; 14'h 54f: x = 16'h4767; 14'h 550: x = 16'h4764; 14'h 551: x = 16'h4762; 14'h 552: x = 16'h475f; 14'h 553: x = 16'h475c; 14'h 554: x = 16'h475a; 14'h 555: x = 16'h4757; 14'h 556: x = 16'h4754; 14'h 557: x = 16'h4752; 14'h 558: x = 16'h474f; 14'h 559: x = 16'h474c; 14'h 55a: x = 16'h4749; 14'h 55b: x = 16'h4747; 14'h 55c: x = 16'h4744; 14'h 55d: x = 16'h4741; 14'h 55e: x = 16'h473f; 14'h 55f: x = 16'h473c; 14'h 560: x = 16'h4739; 14'h 561: x = 16'h4737; 14'h 562: x = 16'h4734; 14'h 563: x = 16'h4731; 14'h 564: x = 16'h472f; 14'h 565: x = 16'h472c; 14'h 566: x = 16'h4729; 14'h 567: x = 16'h4727; 14'h 568: x = 16'h4724; 14'h 569: x = 16'h4721; 14'h 56a: x = 16'h471f; 14'h 56b: x = 16'h471c; 14'h 56c: x = 16'h4719; 14'h 56d: x = 16'h4717; 14'h 56e: x = 16'h4714; 14'h 56f: x = 16'h4711; 14'h 570: x = 16'h470f; 14'h 571: x = 16'h470c; 14'h 572: x = 16'h4709; 14'h 573: x = 16'h4707; 14'h 574: x = 16'h4704; 14'h 575: x = 16'h4702; 14'h 576: x = 16'h46ff; 14'h 577: x = 16'h46fc; 14'h 578: x = 16'h46fa; 14'h 579: x = 16'h46f7; 14'h 57a: x = 16'h46f4; 14'h 57b: x = 16'h46f2; 14'h 57c: x = 16'h46ef; 14'h 57d: x = 16'h46ec; 14'h 57e: x = 16'h46ea; 14'h 57f: x = 16'h46e7; 14'h 580: x = 16'h46e5; 14'h 581: x = 16'h46e2; 14'h 582: x = 16'h46df; 14'h 583: x = 16'h46dd; 14'h 584: x = 16'h46da; 14'h 585: x = 16'h46d7; 14'h 586: x = 16'h46d5; 14'h 587: x = 16'h46d2; 14'h 588: x = 16'h46d0; 14'h 589: x = 16'h46cd; 14'h 58a: x = 16'h46ca; 14'h 58b: x = 16'h46c8; 14'h 58c: x = 16'h46c5; 14'h 58d: x = 16'h46c3; 14'h 58e: x = 16'h46c0; 14'h 58f: x = 16'h46bd; 14'h 590: x = 16'h46bb; 14'h 591: x = 16'h46b8; 14'h 592: x = 16'h46b6; 14'h 593: x = 16'h46b3; 14'h 594: x = 16'h46b0; 14'h 595: x = 16'h46ae; 14'h 596: x = 16'h46ab; 14'h 597: x = 16'h46a9; 14'h 598: x = 16'h46a6; 14'h 599: x = 16'h46a3; 14'h 59a: x = 16'h46a1; 14'h 59b: x = 16'h469e; 14'h 59c: x = 16'h469c; 14'h 59d: x = 16'h4699; 14'h 59e: x = 16'h4696; 14'h 59f: x = 16'h4694; 14'h 5a0: x = 16'h4691; 14'h 5a1: x = 16'h468f; 14'h 5a2: x = 16'h468c; 14'h 5a3: x = 16'h468a; 14'h 5a4: x = 16'h4687; 14'h 5a5: x = 16'h4684; 14'h 5a6: x = 16'h4682; 14'h 5a7: x = 16'h467f; 14'h 5a8: x = 16'h467d; 14'h 5a9: x = 16'h467a; 14'h 5aa: x = 16'h4678; 14'h 5ab: x = 16'h4675; 14'h 5ac: x = 16'h4672; 14'h 5ad: x = 16'h4670; 14'h 5ae: x = 16'h466d; 14'h 5af: x = 16'h466b; 14'h 5b0: x = 16'h4668; 14'h 5b1: x = 16'h4666; 14'h 5b2: x = 16'h4663; 14'h 5b3: x = 16'h4661; 14'h 5b4: x = 16'h465e; 14'h 5b5: x = 16'h465b; 14'h 5b6: x = 16'h4659; 14'h 5b7: x = 16'h4656; 14'h 5b8: x = 16'h4654; 14'h 5b9: x = 16'h4651; 14'h 5ba: x = 16'h464f; 14'h 5bb: x = 16'h464c; 14'h 5bc: x = 16'h464a; 14'h 5bd: x = 16'h4647; 14'h 5be: x = 16'h4645; 14'h 5bf: x = 16'h4642; 14'h 5c0: x = 16'h463f; 14'h 5c1: x = 16'h463d; 14'h 5c2: x = 16'h463a; 14'h 5c3: x = 16'h4638; 14'h 5c4: x = 16'h4635; 14'h 5c5: x = 16'h4633; 14'h 5c6: x = 16'h4630; 14'h 5c7: x = 16'h462e; 14'h 5c8: x = 16'h462b; 14'h 5c9: x = 16'h4629; 14'h 5ca: x = 16'h4626; 14'h 5cb: x = 16'h4624; 14'h 5cc: x = 16'h4621; 14'h 5cd: x = 16'h461f; 14'h 5ce: x = 16'h461c; 14'h 5cf: x = 16'h461a; 14'h 5d0: x = 16'h4617; 14'h 5d1: x = 16'h4615; 14'h 5d2: x = 16'h4612; 14'h 5d3: x = 16'h4610; 14'h 5d4: x = 16'h460d; 14'h 5d5: x = 16'h460b; 14'h 5d6: x = 16'h4608; 14'h 5d7: x = 16'h4605; 14'h 5d8: x = 16'h4603; 14'h 5d9: x = 16'h4600; 14'h 5da: x = 16'h45fe; 14'h 5db: x = 16'h45fb; 14'h 5dc: x = 16'h45f9; 14'h 5dd: x = 16'h45f6; 14'h 5de: x = 16'h45f4; 14'h 5df: x = 16'h45f2; 14'h 5e0: x = 16'h45ef; 14'h 5e1: x = 16'h45ed; 14'h 5e2: x = 16'h45ea; 14'h 5e3: x = 16'h45e8; 14'h 5e4: x = 16'h45e5; 14'h 5e5: x = 16'h45e3; 14'h 5e6: x = 16'h45e0; 14'h 5e7: x = 16'h45de; 14'h 5e8: x = 16'h45db; 14'h 5e9: x = 16'h45d9; 14'h 5ea: x = 16'h45d6; 14'h 5eb: x = 16'h45d4; 14'h 5ec: x = 16'h45d1; 14'h 5ed: x = 16'h45cf; 14'h 5ee: x = 16'h45cc; 14'h 5ef: x = 16'h45ca; 14'h 5f0: x = 16'h45c7; 14'h 5f1: x = 16'h45c5; 14'h 5f2: x = 16'h45c2; 14'h 5f3: x = 16'h45c0; 14'h 5f4: x = 16'h45bd; 14'h 5f5: x = 16'h45bb; 14'h 5f6: x = 16'h45b8; 14'h 5f7: x = 16'h45b6; 14'h 5f8: x = 16'h45b4; 14'h 5f9: x = 16'h45b1; 14'h 5fa: x = 16'h45af; 14'h 5fb: x = 16'h45ac; 14'h 5fc: x = 16'h45aa; 14'h 5fd: x = 16'h45a7; 14'h 5fe: x = 16'h45a5; 14'h 5ff: x = 16'h45a2; 14'h 600: x = 16'h45a0; 14'h 601: x = 16'h459d; 14'h 602: x = 16'h459b; 14'h 603: x = 16'h4599; 14'h 604: x = 16'h4596; 14'h 605: x = 16'h4594; 14'h 606: x = 16'h4591; 14'h 607: x = 16'h458f; 14'h 608: x = 16'h458c; 14'h 609: x = 16'h458a; 14'h 60a: x = 16'h4587; 14'h 60b: x = 16'h4585; 14'h 60c: x = 16'h4583; 14'h 60d: x = 16'h4580; 14'h 60e: x = 16'h457e; 14'h 60f: x = 16'h457b; 14'h 610: x = 16'h4579; 14'h 611: x = 16'h4576; 14'h 612: x = 16'h4574; 14'h 613: x = 16'h4572; 14'h 614: x = 16'h456f; 14'h 615: x = 16'h456d; 14'h 616: x = 16'h456a; 14'h 617: x = 16'h4568; 14'h 618: x = 16'h4565; 14'h 619: x = 16'h4563; 14'h 61a: x = 16'h4561; 14'h 61b: x = 16'h455e; 14'h 61c: x = 16'h455c; 14'h 61d: x = 16'h4559; 14'h 61e: x = 16'h4557; 14'h 61f: x = 16'h4555; 14'h 620: x = 16'h4552; 14'h 621: x = 16'h4550; 14'h 622: x = 16'h454d; 14'h 623: x = 16'h454b; 14'h 624: x = 16'h4548; 14'h 625: x = 16'h4546; 14'h 626: x = 16'h4544; 14'h 627: x = 16'h4541; 14'h 628: x = 16'h453f; 14'h 629: x = 16'h453c; 14'h 62a: x = 16'h453a; 14'h 62b: x = 16'h4538; 14'h 62c: x = 16'h4535; 14'h 62d: x = 16'h4533; 14'h 62e: x = 16'h4530; 14'h 62f: x = 16'h452e; 14'h 630: x = 16'h452c; 14'h 631: x = 16'h4529; 14'h 632: x = 16'h4527; 14'h 633: x = 16'h4525; 14'h 634: x = 16'h4522; 14'h 635: x = 16'h4520; 14'h 636: x = 16'h451d; 14'h 637: x = 16'h451b; 14'h 638: x = 16'h4519; 14'h 639: x = 16'h4516; 14'h 63a: x = 16'h4514; 14'h 63b: x = 16'h4511; 14'h 63c: x = 16'h450f; 14'h 63d: x = 16'h450d; 14'h 63e: x = 16'h450a; 14'h 63f: x = 16'h4508; 14'h 640: x = 16'h4506; 14'h 641: x = 16'h4503; 14'h 642: x = 16'h4501; 14'h 643: x = 16'h44fe; 14'h 644: x = 16'h44fc; 14'h 645: x = 16'h44fa; 14'h 646: x = 16'h44f7; 14'h 647: x = 16'h44f5; 14'h 648: x = 16'h44f3; 14'h 649: x = 16'h44f0; 14'h 64a: x = 16'h44ee; 14'h 64b: x = 16'h44ec; 14'h 64c: x = 16'h44e9; 14'h 64d: x = 16'h44e7; 14'h 64e: x = 16'h44e4; 14'h 64f: x = 16'h44e2; 14'h 650: x = 16'h44e0; 14'h 651: x = 16'h44dd; 14'h 652: x = 16'h44db; 14'h 653: x = 16'h44d9; 14'h 654: x = 16'h44d6; 14'h 655: x = 16'h44d4; 14'h 656: x = 16'h44d2; 14'h 657: x = 16'h44cf; 14'h 658: x = 16'h44cd; 14'h 659: x = 16'h44cb; 14'h 65a: x = 16'h44c8; 14'h 65b: x = 16'h44c6; 14'h 65c: x = 16'h44c4; 14'h 65d: x = 16'h44c1; 14'h 65e: x = 16'h44bf; 14'h 65f: x = 16'h44bd; 14'h 660: x = 16'h44ba; 14'h 661: x = 16'h44b8; 14'h 662: x = 16'h44b6; 14'h 663: x = 16'h44b3; 14'h 664: x = 16'h44b1; 14'h 665: x = 16'h44af; 14'h 666: x = 16'h44ac; 14'h 667: x = 16'h44aa; 14'h 668: x = 16'h44a8; 14'h 669: x = 16'h44a5; 14'h 66a: x = 16'h44a3; 14'h 66b: x = 16'h44a1; 14'h 66c: x = 16'h449e; 14'h 66d: x = 16'h449c; 14'h 66e: x = 16'h449a; 14'h 66f: x = 16'h4497; 14'h 670: x = 16'h4495; 14'h 671: x = 16'h4493; 14'h 672: x = 16'h4490; 14'h 673: x = 16'h448e; 14'h 674: x = 16'h448c; 14'h 675: x = 16'h4489; 14'h 676: x = 16'h4487; 14'h 677: x = 16'h4485; 14'h 678: x = 16'h4482; 14'h 679: x = 16'h4480; 14'h 67a: x = 16'h447e; 14'h 67b: x = 16'h447b; 14'h 67c: x = 16'h4479; 14'h 67d: x = 16'h4477; 14'h 67e: x = 16'h4475; 14'h 67f: x = 16'h4472; 14'h 680: x = 16'h4470; 14'h 681: x = 16'h446e; 14'h 682: x = 16'h446b; 14'h 683: x = 16'h4469; 14'h 684: x = 16'h4467; 14'h 685: x = 16'h4464; 14'h 686: x = 16'h4462; 14'h 687: x = 16'h4460; 14'h 688: x = 16'h445e; 14'h 689: x = 16'h445b; 14'h 68a: x = 16'h4459; 14'h 68b: x = 16'h4457; 14'h 68c: x = 16'h4454; 14'h 68d: x = 16'h4452; 14'h 68e: x = 16'h4450; 14'h 68f: x = 16'h444e; 14'h 690: x = 16'h444b; 14'h 691: x = 16'h4449; 14'h 692: x = 16'h4447; 14'h 693: x = 16'h4444; 14'h 694: x = 16'h4442; 14'h 695: x = 16'h4440; 14'h 696: x = 16'h443e; 14'h 697: x = 16'h443b; 14'h 698: x = 16'h4439; 14'h 699: x = 16'h4437; 14'h 69a: x = 16'h4434; 14'h 69b: x = 16'h4432; 14'h 69c: x = 16'h4430; 14'h 69d: x = 16'h442e; 14'h 69e: x = 16'h442b; 14'h 69f: x = 16'h4429; 14'h 6a0: x = 16'h4427; 14'h 6a1: x = 16'h4425; 14'h 6a2: x = 16'h4422; 14'h 6a3: x = 16'h4420; 14'h 6a4: x = 16'h441e; 14'h 6a5: x = 16'h441c; 14'h 6a6: x = 16'h4419; 14'h 6a7: x = 16'h4417; 14'h 6a8: x = 16'h4415; 14'h 6a9: x = 16'h4412; 14'h 6aa: x = 16'h4410; 14'h 6ab: x = 16'h440e; 14'h 6ac: x = 16'h440c; 14'h 6ad: x = 16'h4409; 14'h 6ae: x = 16'h4407; 14'h 6af: x = 16'h4405; 14'h 6b0: x = 16'h4403; 14'h 6b1: x = 16'h4400; 14'h 6b2: x = 16'h43fe; 14'h 6b3: x = 16'h43fc; 14'h 6b4: x = 16'h43fa; 14'h 6b5: x = 16'h43f7; 14'h 6b6: x = 16'h43f5; 14'h 6b7: x = 16'h43f3; 14'h 6b8: x = 16'h43f1; 14'h 6b9: x = 16'h43ee; 14'h 6ba: x = 16'h43ec; 14'h 6bb: x = 16'h43ea; 14'h 6bc: x = 16'h43e8; 14'h 6bd: x = 16'h43e6; 14'h 6be: x = 16'h43e3; 14'h 6bf: x = 16'h43e1; 14'h 6c0: x = 16'h43df; 14'h 6c1: x = 16'h43dd; 14'h 6c2: x = 16'h43da; 14'h 6c3: x = 16'h43d8; 14'h 6c4: x = 16'h43d6; 14'h 6c5: x = 16'h43d4; 14'h 6c6: x = 16'h43d1; 14'h 6c7: x = 16'h43cf; 14'h 6c8: x = 16'h43cd; 14'h 6c9: x = 16'h43cb; 14'h 6ca: x = 16'h43c9; 14'h 6cb: x = 16'h43c6; 14'h 6cc: x = 16'h43c4; 14'h 6cd: x = 16'h43c2; 14'h 6ce: x = 16'h43c0; 14'h 6cf: x = 16'h43bd; 14'h 6d0: x = 16'h43bb; 14'h 6d1: x = 16'h43b9; 14'h 6d2: x = 16'h43b7; 14'h 6d3: x = 16'h43b5; 14'h 6d4: x = 16'h43b2; 14'h 6d5: x = 16'h43b0; 14'h 6d6: x = 16'h43ae; 14'h 6d7: x = 16'h43ac; 14'h 6d8: x = 16'h43a9; 14'h 6d9: x = 16'h43a7; 14'h 6da: x = 16'h43a5; 14'h 6db: x = 16'h43a3; 14'h 6dc: x = 16'h43a1; 14'h 6dd: x = 16'h439e; 14'h 6de: x = 16'h439c; 14'h 6df: x = 16'h439a; 14'h 6e0: x = 16'h4398; 14'h 6e1: x = 16'h4396; 14'h 6e2: x = 16'h4393; 14'h 6e3: x = 16'h4391; 14'h 6e4: x = 16'h438f; 14'h 6e5: x = 16'h438d; 14'h 6e6: x = 16'h438b; 14'h 6e7: x = 16'h4388; 14'h 6e8: x = 16'h4386; 14'h 6e9: x = 16'h4384; 14'h 6ea: x = 16'h4382; 14'h 6eb: x = 16'h4380; 14'h 6ec: x = 16'h437d; 14'h 6ed: x = 16'h437b; 14'h 6ee: x = 16'h4379; 14'h 6ef: x = 16'h4377; 14'h 6f0: x = 16'h4375; 14'h 6f1: x = 16'h4372; 14'h 6f2: x = 16'h4370; 14'h 6f3: x = 16'h436e; 14'h 6f4: x = 16'h436c; 14'h 6f5: x = 16'h436a; 14'h 6f6: x = 16'h4368; 14'h 6f7: x = 16'h4365; 14'h 6f8: x = 16'h4363; 14'h 6f9: x = 16'h4361; 14'h 6fa: x = 16'h435f; 14'h 6fb: x = 16'h435d; 14'h 6fc: x = 16'h435a; 14'h 6fd: x = 16'h4358; 14'h 6fe: x = 16'h4356; 14'h 6ff: x = 16'h4354; 14'h 700: x = 16'h4352; 14'h 701: x = 16'h4350; 14'h 702: x = 16'h434d; 14'h 703: x = 16'h434b; 14'h 704: x = 16'h4349; 14'h 705: x = 16'h4347; 14'h 706: x = 16'h4345; 14'h 707: x = 16'h4343; 14'h 708: x = 16'h4340; 14'h 709: x = 16'h433e; 14'h 70a: x = 16'h433c; 14'h 70b: x = 16'h433a; 14'h 70c: x = 16'h4338; 14'h 70d: x = 16'h4336; 14'h 70e: x = 16'h4333; 14'h 70f: x = 16'h4331; 14'h 710: x = 16'h432f; 14'h 711: x = 16'h432d; 14'h 712: x = 16'h432b; 14'h 713: x = 16'h4329; 14'h 714: x = 16'h4327; 14'h 715: x = 16'h4324; 14'h 716: x = 16'h4322; 14'h 717: x = 16'h4320; 14'h 718: x = 16'h431e; 14'h 719: x = 16'h431c; 14'h 71a: x = 16'h431a; 14'h 71b: x = 16'h4317; 14'h 71c: x = 16'h4315; 14'h 71d: x = 16'h4313; 14'h 71e: x = 16'h4311; 14'h 71f: x = 16'h430f; 14'h 720: x = 16'h430d; 14'h 721: x = 16'h430b; 14'h 722: x = 16'h4308; 14'h 723: x = 16'h4306; 14'h 724: x = 16'h4304; 14'h 725: x = 16'h4302; 14'h 726: x = 16'h4300; 14'h 727: x = 16'h42fe; 14'h 728: x = 16'h42fc; 14'h 729: x = 16'h42f9; 14'h 72a: x = 16'h42f7; 14'h 72b: x = 16'h42f5; 14'h 72c: x = 16'h42f3; 14'h 72d: x = 16'h42f1; 14'h 72e: x = 16'h42ef; 14'h 72f: x = 16'h42ed; 14'h 730: x = 16'h42eb; 14'h 731: x = 16'h42e8; 14'h 732: x = 16'h42e6; 14'h 733: x = 16'h42e4; 14'h 734: x = 16'h42e2; 14'h 735: x = 16'h42e0; 14'h 736: x = 16'h42de; 14'h 737: x = 16'h42dc; 14'h 738: x = 16'h42da; 14'h 739: x = 16'h42d7; 14'h 73a: x = 16'h42d5; 14'h 73b: x = 16'h42d3; 14'h 73c: x = 16'h42d1; 14'h 73d: x = 16'h42cf; 14'h 73e: x = 16'h42cd; 14'h 73f: x = 16'h42cb; 14'h 740: x = 16'h42c9; 14'h 741: x = 16'h42c6; 14'h 742: x = 16'h42c4; 14'h 743: x = 16'h42c2; 14'h 744: x = 16'h42c0; 14'h 745: x = 16'h42be; 14'h 746: x = 16'h42bc; 14'h 747: x = 16'h42ba; 14'h 748: x = 16'h42b8; 14'h 749: x = 16'h42b6; 14'h 74a: x = 16'h42b3; 14'h 74b: x = 16'h42b1; 14'h 74c: x = 16'h42af; 14'h 74d: x = 16'h42ad; 14'h 74e: x = 16'h42ab; 14'h 74f: x = 16'h42a9; 14'h 750: x = 16'h42a7; 14'h 751: x = 16'h42a5; 14'h 752: x = 16'h42a3; 14'h 753: x = 16'h42a1; 14'h 754: x = 16'h429e; 14'h 755: x = 16'h429c; 14'h 756: x = 16'h429a; 14'h 757: x = 16'h4298; 14'h 758: x = 16'h4296; 14'h 759: x = 16'h4294; 14'h 75a: x = 16'h4292; 14'h 75b: x = 16'h4290; 14'h 75c: x = 16'h428e; 14'h 75d: x = 16'h428c; 14'h 75e: x = 16'h428a; 14'h 75f: x = 16'h4287; 14'h 760: x = 16'h4285; 14'h 761: x = 16'h4283; 14'h 762: x = 16'h4281; 14'h 763: x = 16'h427f; 14'h 764: x = 16'h427d; 14'h 765: x = 16'h427b; 14'h 766: x = 16'h4279; 14'h 767: x = 16'h4277; 14'h 768: x = 16'h4275; 14'h 769: x = 16'h4273; 14'h 76a: x = 16'h4271; 14'h 76b: x = 16'h426e; 14'h 76c: x = 16'h426c; 14'h 76d: x = 16'h426a; 14'h 76e: x = 16'h4268; 14'h 76f: x = 16'h4266; 14'h 770: x = 16'h4264; 14'h 771: x = 16'h4262; 14'h 772: x = 16'h4260; 14'h 773: x = 16'h425e; 14'h 774: x = 16'h425c; 14'h 775: x = 16'h425a; 14'h 776: x = 16'h4258; 14'h 777: x = 16'h4256; 14'h 778: x = 16'h4254; 14'h 779: x = 16'h4251; 14'h 77a: x = 16'h424f; 14'h 77b: x = 16'h424d; 14'h 77c: x = 16'h424b; 14'h 77d: x = 16'h4249; 14'h 77e: x = 16'h4247; 14'h 77f: x = 16'h4245; 14'h 780: x = 16'h4243; 14'h 781: x = 16'h4241; 14'h 782: x = 16'h423f; 14'h 783: x = 16'h423d; 14'h 784: x = 16'h423b; 14'h 785: x = 16'h4239; 14'h 786: x = 16'h4237; 14'h 787: x = 16'h4235; 14'h 788: x = 16'h4233; 14'h 789: x = 16'h4230; 14'h 78a: x = 16'h422e; 14'h 78b: x = 16'h422c; 14'h 78c: x = 16'h422a; 14'h 78d: x = 16'h4228; 14'h 78e: x = 16'h4226; 14'h 78f: x = 16'h4224; 14'h 790: x = 16'h4222; 14'h 791: x = 16'h4220; 14'h 792: x = 16'h421e; 14'h 793: x = 16'h421c; 14'h 794: x = 16'h421a; 14'h 795: x = 16'h4218; 14'h 796: x = 16'h4216; 14'h 797: x = 16'h4214; 14'h 798: x = 16'h4212; 14'h 799: x = 16'h4210; 14'h 79a: x = 16'h420e; 14'h 79b: x = 16'h420c; 14'h 79c: x = 16'h420a; 14'h 79d: x = 16'h4208; 14'h 79e: x = 16'h4206; 14'h 79f: x = 16'h4204; 14'h 7a0: x = 16'h4201; 14'h 7a1: x = 16'h41ff; 14'h 7a2: x = 16'h41fd; 14'h 7a3: x = 16'h41fb; 14'h 7a4: x = 16'h41f9; 14'h 7a5: x = 16'h41f7; 14'h 7a6: x = 16'h41f5; 14'h 7a7: x = 16'h41f3; 14'h 7a8: x = 16'h41f1; 14'h 7a9: x = 16'h41ef; 14'h 7aa: x = 16'h41ed; 14'h 7ab: x = 16'h41eb; 14'h 7ac: x = 16'h41e9; 14'h 7ad: x = 16'h41e7; 14'h 7ae: x = 16'h41e5; 14'h 7af: x = 16'h41e3; 14'h 7b0: x = 16'h41e1; 14'h 7b1: x = 16'h41df; 14'h 7b2: x = 16'h41dd; 14'h 7b3: x = 16'h41db; 14'h 7b4: x = 16'h41d9; 14'h 7b5: x = 16'h41d7; 14'h 7b6: x = 16'h41d5; 14'h 7b7: x = 16'h41d3; 14'h 7b8: x = 16'h41d1; 14'h 7b9: x = 16'h41cf; 14'h 7ba: x = 16'h41cd; 14'h 7bb: x = 16'h41cb; 14'h 7bc: x = 16'h41c9; 14'h 7bd: x = 16'h41c7; 14'h 7be: x = 16'h41c5; 14'h 7bf: x = 16'h41c3; 14'h 7c0: x = 16'h41c1; 14'h 7c1: x = 16'h41bf; 14'h 7c2: x = 16'h41bd; 14'h 7c3: x = 16'h41bb; 14'h 7c4: x = 16'h41b9; 14'h 7c5: x = 16'h41b7; 14'h 7c6: x = 16'h41b5; 14'h 7c7: x = 16'h41b3; 14'h 7c8: x = 16'h41b1; 14'h 7c9: x = 16'h41af; 14'h 7ca: x = 16'h41ad; 14'h 7cb: x = 16'h41ab; 14'h 7cc: x = 16'h41a9; 14'h 7cd: x = 16'h41a7; 14'h 7ce: x = 16'h41a5; 14'h 7cf: x = 16'h41a3; 14'h 7d0: x = 16'h41a1; 14'h 7d1: x = 16'h419f; 14'h 7d2: x = 16'h419d; 14'h 7d3: x = 16'h419b; 14'h 7d4: x = 16'h4199; 14'h 7d5: x = 16'h4197; 14'h 7d6: x = 16'h4195; 14'h 7d7: x = 16'h4193; 14'h 7d8: x = 16'h4191; 14'h 7d9: x = 16'h418f; 14'h 7da: x = 16'h418d; 14'h 7db: x = 16'h418b; 14'h 7dc: x = 16'h4189; 14'h 7dd: x = 16'h4187; 14'h 7de: x = 16'h4185; 14'h 7df: x = 16'h4183; 14'h 7e0: x = 16'h4181; 14'h 7e1: x = 16'h417f; 14'h 7e2: x = 16'h417d; 14'h 7e3: x = 16'h417b; 14'h 7e4: x = 16'h4179; 14'h 7e5: x = 16'h4177; 14'h 7e6: x = 16'h4175; 14'h 7e7: x = 16'h4173; 14'h 7e8: x = 16'h4171; 14'h 7e9: x = 16'h416f; 14'h 7ea: x = 16'h416d; 14'h 7eb: x = 16'h416b; 14'h 7ec: x = 16'h4169; 14'h 7ed: x = 16'h4167; 14'h 7ee: x = 16'h4165; 14'h 7ef: x = 16'h4163; 14'h 7f0: x = 16'h4161; 14'h 7f1: x = 16'h415f; 14'h 7f2: x = 16'h415d; 14'h 7f3: x = 16'h415b; 14'h 7f4: x = 16'h4159; 14'h 7f5: x = 16'h4157; 14'h 7f6: x = 16'h4155; 14'h 7f7: x = 16'h4153; 14'h 7f8: x = 16'h4151; 14'h 7f9: x = 16'h414f; 14'h 7fa: x = 16'h414e; 14'h 7fb: x = 16'h414c; 14'h 7fc: x = 16'h414a; 14'h 7fd: x = 16'h4148; 14'h 7fe: x = 16'h4146; 14'h 7ff: x = 16'h4144; 14'h 800: x = 16'h4142; 14'h 801: x = 16'h4140; 14'h 802: x = 16'h413e; 14'h 803: x = 16'h413c; 14'h 804: x = 16'h413a; 14'h 805: x = 16'h4138; 14'h 806: x = 16'h4136; 14'h 807: x = 16'h4134; 14'h 808: x = 16'h4132; 14'h 809: x = 16'h4130; 14'h 80a: x = 16'h412e; 14'h 80b: x = 16'h412c; 14'h 80c: x = 16'h412a; 14'h 80d: x = 16'h4128; 14'h 80e: x = 16'h4126; 14'h 80f: x = 16'h4124; 14'h 810: x = 16'h4122; 14'h 811: x = 16'h4120; 14'h 812: x = 16'h411f; 14'h 813: x = 16'h411d; 14'h 814: x = 16'h411b; 14'h 815: x = 16'h4119; 14'h 816: x = 16'h4117; 14'h 817: x = 16'h4115; 14'h 818: x = 16'h4113; 14'h 819: x = 16'h4111; 14'h 81a: x = 16'h410f; 14'h 81b: x = 16'h410d; 14'h 81c: x = 16'h410b; 14'h 81d: x = 16'h4109; 14'h 81e: x = 16'h4107; 14'h 81f: x = 16'h4105; 14'h 820: x = 16'h4103; 14'h 821: x = 16'h4101; 14'h 822: x = 16'h40ff; 14'h 823: x = 16'h40fe; 14'h 824: x = 16'h40fc; 14'h 825: x = 16'h40fa; 14'h 826: x = 16'h40f8; 14'h 827: x = 16'h40f6; 14'h 828: x = 16'h40f4; 14'h 829: x = 16'h40f2; 14'h 82a: x = 16'h40f0; 14'h 82b: x = 16'h40ee; 14'h 82c: x = 16'h40ec; 14'h 82d: x = 16'h40ea; 14'h 82e: x = 16'h40e8; 14'h 82f: x = 16'h40e6; 14'h 830: x = 16'h40e4; 14'h 831: x = 16'h40e2; 14'h 832: x = 16'h40e1; 14'h 833: x = 16'h40df; 14'h 834: x = 16'h40dd; 14'h 835: x = 16'h40db; 14'h 836: x = 16'h40d9; 14'h 837: x = 16'h40d7; 14'h 838: x = 16'h40d5; 14'h 839: x = 16'h40d3; 14'h 83a: x = 16'h40d1; 14'h 83b: x = 16'h40cf; 14'h 83c: x = 16'h40cd; 14'h 83d: x = 16'h40cb; 14'h 83e: x = 16'h40c9; 14'h 83f: x = 16'h40c8; 14'h 840: x = 16'h40c6; 14'h 841: x = 16'h40c4; 14'h 842: x = 16'h40c2; 14'h 843: x = 16'h40c0; 14'h 844: x = 16'h40be; 14'h 845: x = 16'h40bc; 14'h 846: x = 16'h40ba; 14'h 847: x = 16'h40b8; 14'h 848: x = 16'h40b6; 14'h 849: x = 16'h40b4; 14'h 84a: x = 16'h40b3; 14'h 84b: x = 16'h40b1; 14'h 84c: x = 16'h40af; 14'h 84d: x = 16'h40ad; 14'h 84e: x = 16'h40ab; 14'h 84f: x = 16'h40a9; 14'h 850: x = 16'h40a7; 14'h 851: x = 16'h40a5; 14'h 852: x = 16'h40a3; 14'h 853: x = 16'h40a1; 14'h 854: x = 16'h409f; 14'h 855: x = 16'h409e; 14'h 856: x = 16'h409c; 14'h 857: x = 16'h409a; 14'h 858: x = 16'h4098; 14'h 859: x = 16'h4096; 14'h 85a: x = 16'h4094; 14'h 85b: x = 16'h4092; 14'h 85c: x = 16'h4090; 14'h 85d: x = 16'h408e; 14'h 85e: x = 16'h408c; 14'h 85f: x = 16'h408b; 14'h 860: x = 16'h4089; 14'h 861: x = 16'h4087; 14'h 862: x = 16'h4085; 14'h 863: x = 16'h4083; 14'h 864: x = 16'h4081; 14'h 865: x = 16'h407f; 14'h 866: x = 16'h407d; 14'h 867: x = 16'h407b; 14'h 868: x = 16'h407a; 14'h 869: x = 16'h4078; 14'h 86a: x = 16'h4076; 14'h 86b: x = 16'h4074; 14'h 86c: x = 16'h4072; 14'h 86d: x = 16'h4070; 14'h 86e: x = 16'h406e; 14'h 86f: x = 16'h406c; 14'h 870: x = 16'h406a; 14'h 871: x = 16'h4069; 14'h 872: x = 16'h4067; 14'h 873: x = 16'h4065; 14'h 874: x = 16'h4063; 14'h 875: x = 16'h4061; 14'h 876: x = 16'h405f; 14'h 877: x = 16'h405d; 14'h 878: x = 16'h405b; 14'h 879: x = 16'h405a; 14'h 87a: x = 16'h4058; 14'h 87b: x = 16'h4056; 14'h 87c: x = 16'h4054; 14'h 87d: x = 16'h4052; 14'h 87e: x = 16'h4050; 14'h 87f: x = 16'h404e; 14'h 880: x = 16'h404c; 14'h 881: x = 16'h404b; 14'h 882: x = 16'h4049; 14'h 883: x = 16'h4047; 14'h 884: x = 16'h4045; 14'h 885: x = 16'h4043; 14'h 886: x = 16'h4041; 14'h 887: x = 16'h403f; 14'h 888: x = 16'h403d; 14'h 889: x = 16'h403c; 14'h 88a: x = 16'h403a; 14'h 88b: x = 16'h4038; 14'h 88c: x = 16'h4036; 14'h 88d: x = 16'h4034; 14'h 88e: x = 16'h4032; 14'h 88f: x = 16'h4030; 14'h 890: x = 16'h402e; 14'h 891: x = 16'h402d; 14'h 892: x = 16'h402b; 14'h 893: x = 16'h4029; 14'h 894: x = 16'h4027; 14'h 895: x = 16'h4025; 14'h 896: x = 16'h4023; 14'h 897: x = 16'h4021; 14'h 898: x = 16'h4020; 14'h 899: x = 16'h401e; 14'h 89a: x = 16'h401c; 14'h 89b: x = 16'h401a; 14'h 89c: x = 16'h4018; 14'h 89d: x = 16'h4016; 14'h 89e: x = 16'h4014; 14'h 89f: x = 16'h4013; 14'h 8a0: x = 16'h4011; 14'h 8a1: x = 16'h400f; 14'h 8a2: x = 16'h400d; 14'h 8a3: x = 16'h400b; 14'h 8a4: x = 16'h4009; 14'h 8a5: x = 16'h4008; 14'h 8a6: x = 16'h4006; 14'h 8a7: x = 16'h4004; 14'h 8a8: x = 16'h4002; 14'h 8a9: x = 16'h4000; 14'h 8aa: x = 16'h3ffe; 14'h 8ab: x = 16'h3ffc; 14'h 8ac: x = 16'h3ffb; 14'h 8ad: x = 16'h3ff9; 14'h 8ae: x = 16'h3ff7; 14'h 8af: x = 16'h3ff5; 14'h 8b0: x = 16'h3ff3; 14'h 8b1: x = 16'h3ff1; 14'h 8b2: x = 16'h3ff0; 14'h 8b3: x = 16'h3fee; 14'h 8b4: x = 16'h3fec; 14'h 8b5: x = 16'h3fea; 14'h 8b6: x = 16'h3fe8; 14'h 8b7: x = 16'h3fe6; 14'h 8b8: x = 16'h3fe4; 14'h 8b9: x = 16'h3fe3; 14'h 8ba: x = 16'h3fe1; 14'h 8bb: x = 16'h3fdf; 14'h 8bc: x = 16'h3fdd; 14'h 8bd: x = 16'h3fdb; 14'h 8be: x = 16'h3fd9; 14'h 8bf: x = 16'h3fd8; 14'h 8c0: x = 16'h3fd6; 14'h 8c1: x = 16'h3fd4; 14'h 8c2: x = 16'h3fd2; 14'h 8c3: x = 16'h3fd0; 14'h 8c4: x = 16'h3fce; 14'h 8c5: x = 16'h3fcd; 14'h 8c6: x = 16'h3fcb; 14'h 8c7: x = 16'h3fc9; 14'h 8c8: x = 16'h3fc7; 14'h 8c9: x = 16'h3fc5; 14'h 8ca: x = 16'h3fc3; 14'h 8cb: x = 16'h3fc2; 14'h 8cc: x = 16'h3fc0; 14'h 8cd: x = 16'h3fbe; 14'h 8ce: x = 16'h3fbc; 14'h 8cf: x = 16'h3fba; 14'h 8d0: x = 16'h3fb9; 14'h 8d1: x = 16'h3fb7; 14'h 8d2: x = 16'h3fb5; 14'h 8d3: x = 16'h3fb3; 14'h 8d4: x = 16'h3fb1; 14'h 8d5: x = 16'h3faf; 14'h 8d6: x = 16'h3fae; 14'h 8d7: x = 16'h3fac; 14'h 8d8: x = 16'h3faa; 14'h 8d9: x = 16'h3fa8; 14'h 8da: x = 16'h3fa6; 14'h 8db: x = 16'h3fa5; 14'h 8dc: x = 16'h3fa3; 14'h 8dd: x = 16'h3fa1; 14'h 8de: x = 16'h3f9f; 14'h 8df: x = 16'h3f9d; 14'h 8e0: x = 16'h3f9b; 14'h 8e1: x = 16'h3f9a; 14'h 8e2: x = 16'h3f98; 14'h 8e3: x = 16'h3f96; 14'h 8e4: x = 16'h3f94; 14'h 8e5: x = 16'h3f92; 14'h 8e6: x = 16'h3f91; 14'h 8e7: x = 16'h3f8f; 14'h 8e8: x = 16'h3f8d; 14'h 8e9: x = 16'h3f8b; 14'h 8ea: x = 16'h3f89; 14'h 8eb: x = 16'h3f88; 14'h 8ec: x = 16'h3f86; 14'h 8ed: x = 16'h3f84; 14'h 8ee: x = 16'h3f82; 14'h 8ef: x = 16'h3f80; 14'h 8f0: x = 16'h3f7e; 14'h 8f1: x = 16'h3f7d; 14'h 8f2: x = 16'h3f7b; 14'h 8f3: x = 16'h3f79; 14'h 8f4: x = 16'h3f77; 14'h 8f5: x = 16'h3f75; 14'h 8f6: x = 16'h3f74; 14'h 8f7: x = 16'h3f72; 14'h 8f8: x = 16'h3f70; 14'h 8f9: x = 16'h3f6e; 14'h 8fa: x = 16'h3f6c; 14'h 8fb: x = 16'h3f6b; 14'h 8fc: x = 16'h3f69; 14'h 8fd: x = 16'h3f67; 14'h 8fe: x = 16'h3f65; 14'h 8ff: x = 16'h3f63; 14'h 900: x = 16'h3f62; 14'h 901: x = 16'h3f60; 14'h 902: x = 16'h3f5e; 14'h 903: x = 16'h3f5c; 14'h 904: x = 16'h3f5b; 14'h 905: x = 16'h3f59; 14'h 906: x = 16'h3f57; 14'h 907: x = 16'h3f55; 14'h 908: x = 16'h3f53; 14'h 909: x = 16'h3f52; 14'h 90a: x = 16'h3f50; 14'h 90b: x = 16'h3f4e; 14'h 90c: x = 16'h3f4c; 14'h 90d: x = 16'h3f4a; 14'h 90e: x = 16'h3f49; 14'h 90f: x = 16'h3f47; 14'h 910: x = 16'h3f45; 14'h 911: x = 16'h3f43; 14'h 912: x = 16'h3f41; 14'h 913: x = 16'h3f40; 14'h 914: x = 16'h3f3e; 14'h 915: x = 16'h3f3c; 14'h 916: x = 16'h3f3a; 14'h 917: x = 16'h3f39; 14'h 918: x = 16'h3f37; 14'h 919: x = 16'h3f35; 14'h 91a: x = 16'h3f33; 14'h 91b: x = 16'h3f31; 14'h 91c: x = 16'h3f30; 14'h 91d: x = 16'h3f2e; 14'h 91e: x = 16'h3f2c; 14'h 91f: x = 16'h3f2a; 14'h 920: x = 16'h3f29; 14'h 921: x = 16'h3f27; 14'h 922: x = 16'h3f25; 14'h 923: x = 16'h3f23; 14'h 924: x = 16'h3f21; 14'h 925: x = 16'h3f20; 14'h 926: x = 16'h3f1e; 14'h 927: x = 16'h3f1c; 14'h 928: x = 16'h3f1a; 14'h 929: x = 16'h3f19; 14'h 92a: x = 16'h3f17; 14'h 92b: x = 16'h3f15; 14'h 92c: x = 16'h3f13; 14'h 92d: x = 16'h3f11; 14'h 92e: x = 16'h3f10; 14'h 92f: x = 16'h3f0e; 14'h 930: x = 16'h3f0c; 14'h 931: x = 16'h3f0a; 14'h 932: x = 16'h3f09; 14'h 933: x = 16'h3f07; 14'h 934: x = 16'h3f05; 14'h 935: x = 16'h3f03; 14'h 936: x = 16'h3f02; 14'h 937: x = 16'h3f00; 14'h 938: x = 16'h3efe; 14'h 939: x = 16'h3efc; 14'h 93a: x = 16'h3efb; 14'h 93b: x = 16'h3ef9; 14'h 93c: x = 16'h3ef7; 14'h 93d: x = 16'h3ef5; 14'h 93e: x = 16'h3ef3; 14'h 93f: x = 16'h3ef2; 14'h 940: x = 16'h3ef0; 14'h 941: x = 16'h3eee; 14'h 942: x = 16'h3eec; 14'h 943: x = 16'h3eeb; 14'h 944: x = 16'h3ee9; 14'h 945: x = 16'h3ee7; 14'h 946: x = 16'h3ee5; 14'h 947: x = 16'h3ee4; 14'h 948: x = 16'h3ee2; 14'h 949: x = 16'h3ee0; 14'h 94a: x = 16'h3ede; 14'h 94b: x = 16'h3edd; 14'h 94c: x = 16'h3edb; 14'h 94d: x = 16'h3ed9; 14'h 94e: x = 16'h3ed7; 14'h 94f: x = 16'h3ed6; 14'h 950: x = 16'h3ed4; 14'h 951: x = 16'h3ed2; 14'h 952: x = 16'h3ed0; 14'h 953: x = 16'h3ecf; 14'h 954: x = 16'h3ecd; 14'h 955: x = 16'h3ecb; 14'h 956: x = 16'h3ec9; 14'h 957: x = 16'h3ec8; 14'h 958: x = 16'h3ec6; 14'h 959: x = 16'h3ec4; 14'h 95a: x = 16'h3ec2; 14'h 95b: x = 16'h3ec1; 14'h 95c: x = 16'h3ebf; 14'h 95d: x = 16'h3ebd; 14'h 95e: x = 16'h3ebb; 14'h 95f: x = 16'h3eba; 14'h 960: x = 16'h3eb8; 14'h 961: x = 16'h3eb6; 14'h 962: x = 16'h3eb4; 14'h 963: x = 16'h3eb3; 14'h 964: x = 16'h3eb1; 14'h 965: x = 16'h3eaf; 14'h 966: x = 16'h3eae; 14'h 967: x = 16'h3eac; 14'h 968: x = 16'h3eaa; 14'h 969: x = 16'h3ea8; 14'h 96a: x = 16'h3ea7; 14'h 96b: x = 16'h3ea5; 14'h 96c: x = 16'h3ea3; 14'h 96d: x = 16'h3ea1; 14'h 96e: x = 16'h3ea0; 14'h 96f: x = 16'h3e9e; 14'h 970: x = 16'h3e9c; 14'h 971: x = 16'h3e9a; 14'h 972: x = 16'h3e99; 14'h 973: x = 16'h3e97; 14'h 974: x = 16'h3e95; 14'h 975: x = 16'h3e94; 14'h 976: x = 16'h3e92; 14'h 977: x = 16'h3e90; 14'h 978: x = 16'h3e8e; 14'h 979: x = 16'h3e8d; 14'h 97a: x = 16'h3e8b; 14'h 97b: x = 16'h3e89; 14'h 97c: x = 16'h3e87; 14'h 97d: x = 16'h3e86; 14'h 97e: x = 16'h3e84; 14'h 97f: x = 16'h3e82; 14'h 980: x = 16'h3e81; 14'h 981: x = 16'h3e7f; 14'h 982: x = 16'h3e7d; 14'h 983: x = 16'h3e7b; 14'h 984: x = 16'h3e7a; 14'h 985: x = 16'h3e78; 14'h 986: x = 16'h3e76; 14'h 987: x = 16'h3e74; 14'h 988: x = 16'h3e73; 14'h 989: x = 16'h3e71; 14'h 98a: x = 16'h3e6f; 14'h 98b: x = 16'h3e6e; 14'h 98c: x = 16'h3e6c; 14'h 98d: x = 16'h3e6a; 14'h 98e: x = 16'h3e68; 14'h 98f: x = 16'h3e67; 14'h 990: x = 16'h3e65; 14'h 991: x = 16'h3e63; 14'h 992: x = 16'h3e62; 14'h 993: x = 16'h3e60; 14'h 994: x = 16'h3e5e; 14'h 995: x = 16'h3e5c; 14'h 996: x = 16'h3e5b; 14'h 997: x = 16'h3e59; 14'h 998: x = 16'h3e57; 14'h 999: x = 16'h3e56; 14'h 99a: x = 16'h3e54; 14'h 99b: x = 16'h3e52; 14'h 99c: x = 16'h3e50; 14'h 99d: x = 16'h3e4f; 14'h 99e: x = 16'h3e4d; 14'h 99f: x = 16'h3e4b; 14'h 9a0: x = 16'h3e4a; 14'h 9a1: x = 16'h3e48; 14'h 9a2: x = 16'h3e46; 14'h 9a3: x = 16'h3e44; 14'h 9a4: x = 16'h3e43; 14'h 9a5: x = 16'h3e41; 14'h 9a6: x = 16'h3e3f; 14'h 9a7: x = 16'h3e3e; 14'h 9a8: x = 16'h3e3c; 14'h 9a9: x = 16'h3e3a; 14'h 9aa: x = 16'h3e39; 14'h 9ab: x = 16'h3e37; 14'h 9ac: x = 16'h3e35; 14'h 9ad: x = 16'h3e33; 14'h 9ae: x = 16'h3e32; 14'h 9af: x = 16'h3e30; 14'h 9b0: x = 16'h3e2e; 14'h 9b1: x = 16'h3e2d; 14'h 9b2: x = 16'h3e2b; 14'h 9b3: x = 16'h3e29; 14'h 9b4: x = 16'h3e28; 14'h 9b5: x = 16'h3e26; 14'h 9b6: x = 16'h3e24; 14'h 9b7: x = 16'h3e22; 14'h 9b8: x = 16'h3e21; 14'h 9b9: x = 16'h3e1f; 14'h 9ba: x = 16'h3e1d; 14'h 9bb: x = 16'h3e1c; 14'h 9bc: x = 16'h3e1a; 14'h 9bd: x = 16'h3e18; 14'h 9be: x = 16'h3e17; 14'h 9bf: x = 16'h3e15; 14'h 9c0: x = 16'h3e13; 14'h 9c1: x = 16'h3e12; 14'h 9c2: x = 16'h3e10; 14'h 9c3: x = 16'h3e0e; 14'h 9c4: x = 16'h3e0c; 14'h 9c5: x = 16'h3e0b; 14'h 9c6: x = 16'h3e09; 14'h 9c7: x = 16'h3e07; 14'h 9c8: x = 16'h3e06; 14'h 9c9: x = 16'h3e04; 14'h 9ca: x = 16'h3e02; 14'h 9cb: x = 16'h3e01; 14'h 9cc: x = 16'h3dff; 14'h 9cd: x = 16'h3dfd; 14'h 9ce: x = 16'h3dfc; 14'h 9cf: x = 16'h3dfa; 14'h 9d0: x = 16'h3df8; 14'h 9d1: x = 16'h3df7; 14'h 9d2: x = 16'h3df5; 14'h 9d3: x = 16'h3df3; 14'h 9d4: x = 16'h3df1; 14'h 9d5: x = 16'h3df0; 14'h 9d6: x = 16'h3dee; 14'h 9d7: x = 16'h3dec; 14'h 9d8: x = 16'h3deb; 14'h 9d9: x = 16'h3de9; 14'h 9da: x = 16'h3de7; 14'h 9db: x = 16'h3de6; 14'h 9dc: x = 16'h3de4; 14'h 9dd: x = 16'h3de2; 14'h 9de: x = 16'h3de1; 14'h 9df: x = 16'h3ddf; 14'h 9e0: x = 16'h3ddd; 14'h 9e1: x = 16'h3ddc; 14'h 9e2: x = 16'h3dda; 14'h 9e3: x = 16'h3dd8; 14'h 9e4: x = 16'h3dd7; 14'h 9e5: x = 16'h3dd5; 14'h 9e6: x = 16'h3dd3; 14'h 9e7: x = 16'h3dd2; 14'h 9e8: x = 16'h3dd0; 14'h 9e9: x = 16'h3dce; 14'h 9ea: x = 16'h3dcd; 14'h 9eb: x = 16'h3dcb; 14'h 9ec: x = 16'h3dc9; 14'h 9ed: x = 16'h3dc8; 14'h 9ee: x = 16'h3dc6; 14'h 9ef: x = 16'h3dc4; 14'h 9f0: x = 16'h3dc3; 14'h 9f1: x = 16'h3dc1; 14'h 9f2: x = 16'h3dbf; 14'h 9f3: x = 16'h3dbe; 14'h 9f4: x = 16'h3dbc; 14'h 9f5: x = 16'h3dba; 14'h 9f6: x = 16'h3db9; 14'h 9f7: x = 16'h3db7; 14'h 9f8: x = 16'h3db5; 14'h 9f9: x = 16'h3db4; 14'h 9fa: x = 16'h3db2; 14'h 9fb: x = 16'h3db0; 14'h 9fc: x = 16'h3daf; 14'h 9fd: x = 16'h3dad; 14'h 9fe: x = 16'h3dab; 14'h 9ff: x = 16'h3daa; 14'h a00: x = 16'h3da8; 14'h a01: x = 16'h3da6; 14'h a02: x = 16'h3da5; 14'h a03: x = 16'h3da3; 14'h a04: x = 16'h3da1; 14'h a05: x = 16'h3da0; 14'h a06: x = 16'h3d9e; 14'h a07: x = 16'h3d9c; 14'h a08: x = 16'h3d9b; 14'h a09: x = 16'h3d99; 14'h a0a: x = 16'h3d97; 14'h a0b: x = 16'h3d96; 14'h a0c: x = 16'h3d94; 14'h a0d: x = 16'h3d92; 14'h a0e: x = 16'h3d91; 14'h a0f: x = 16'h3d8f; 14'h a10: x = 16'h3d8d; 14'h a11: x = 16'h3d8c; 14'h a12: x = 16'h3d8a; 14'h a13: x = 16'h3d88; 14'h a14: x = 16'h3d87; 14'h a15: x = 16'h3d85; 14'h a16: x = 16'h3d84; 14'h a17: x = 16'h3d82; 14'h a18: x = 16'h3d80; 14'h a19: x = 16'h3d7f; 14'h a1a: x = 16'h3d7d; 14'h a1b: x = 16'h3d7b; 14'h a1c: x = 16'h3d7a; 14'h a1d: x = 16'h3d78; 14'h a1e: x = 16'h3d76; 14'h a1f: x = 16'h3d75; 14'h a20: x = 16'h3d73; 14'h a21: x = 16'h3d71; 14'h a22: x = 16'h3d70; 14'h a23: x = 16'h3d6e; 14'h a24: x = 16'h3d6c; 14'h a25: x = 16'h3d6b; 14'h a26: x = 16'h3d69; 14'h a27: x = 16'h3d68; 14'h a28: x = 16'h3d66; 14'h a29: x = 16'h3d64; 14'h a2a: x = 16'h3d63; 14'h a2b: x = 16'h3d61; 14'h a2c: x = 16'h3d5f; 14'h a2d: x = 16'h3d5e; 14'h a2e: x = 16'h3d5c; 14'h a2f: x = 16'h3d5a; 14'h a30: x = 16'h3d59; 14'h a31: x = 16'h3d57; 14'h a32: x = 16'h3d55; 14'h a33: x = 16'h3d54; 14'h a34: x = 16'h3d52; 14'h a35: x = 16'h3d51; 14'h a36: x = 16'h3d4f; 14'h a37: x = 16'h3d4d; 14'h a38: x = 16'h3d4c; 14'h a39: x = 16'h3d4a; 14'h a3a: x = 16'h3d48; 14'h a3b: x = 16'h3d47; 14'h a3c: x = 16'h3d45; 14'h a3d: x = 16'h3d43; 14'h a3e: x = 16'h3d42; 14'h a3f: x = 16'h3d40; 14'h a40: x = 16'h3d3f; 14'h a41: x = 16'h3d3d; 14'h a42: x = 16'h3d3b; 14'h a43: x = 16'h3d3a; 14'h a44: x = 16'h3d38; 14'h a45: x = 16'h3d36; 14'h a46: x = 16'h3d35; 14'h a47: x = 16'h3d33; 14'h a48: x = 16'h3d32; 14'h a49: x = 16'h3d30; 14'h a4a: x = 16'h3d2e; 14'h a4b: x = 16'h3d2d; 14'h a4c: x = 16'h3d2b; 14'h a4d: x = 16'h3d29; 14'h a4e: x = 16'h3d28; 14'h a4f: x = 16'h3d26; 14'h a50: x = 16'h3d25; 14'h a51: x = 16'h3d23; 14'h a52: x = 16'h3d21; 14'h a53: x = 16'h3d20; 14'h a54: x = 16'h3d1e; 14'h a55: x = 16'h3d1c; 14'h a56: x = 16'h3d1b; 14'h a57: x = 16'h3d19; 14'h a58: x = 16'h3d18; 14'h a59: x = 16'h3d16; 14'h a5a: x = 16'h3d14; 14'h a5b: x = 16'h3d13; 14'h a5c: x = 16'h3d11; 14'h a5d: x = 16'h3d0f; 14'h a5e: x = 16'h3d0e; 14'h a5f: x = 16'h3d0c; 14'h a60: x = 16'h3d0b; 14'h a61: x = 16'h3d09; 14'h a62: x = 16'h3d07; 14'h a63: x = 16'h3d06; 14'h a64: x = 16'h3d04; 14'h a65: x = 16'h3d03; 14'h a66: x = 16'h3d01; 14'h a67: x = 16'h3cff; 14'h a68: x = 16'h3cfe; 14'h a69: x = 16'h3cfc; 14'h a6a: x = 16'h3cfa; 14'h a6b: x = 16'h3cf9; 14'h a6c: x = 16'h3cf7; 14'h a6d: x = 16'h3cf6; 14'h a6e: x = 16'h3cf4; 14'h a6f: x = 16'h3cf2; 14'h a70: x = 16'h3cf1; 14'h a71: x = 16'h3cef; 14'h a72: x = 16'h3cee; 14'h a73: x = 16'h3cec; 14'h a74: x = 16'h3cea; 14'h a75: x = 16'h3ce9; 14'h a76: x = 16'h3ce7; 14'h a77: x = 16'h3ce6; 14'h a78: x = 16'h3ce4; 14'h a79: x = 16'h3ce2; 14'h a7a: x = 16'h3ce1; 14'h a7b: x = 16'h3cdf; 14'h a7c: x = 16'h3cde; 14'h a7d: x = 16'h3cdc; 14'h a7e: x = 16'h3cda; 14'h a7f: x = 16'h3cd9; 14'h a80: x = 16'h3cd7; 14'h a81: x = 16'h3cd6; 14'h a82: x = 16'h3cd4; 14'h a83: x = 16'h3cd2; 14'h a84: x = 16'h3cd1; 14'h a85: x = 16'h3ccf; 14'h a86: x = 16'h3ccd; 14'h a87: x = 16'h3ccc; 14'h a88: x = 16'h3cca; 14'h a89: x = 16'h3cc9; 14'h a8a: x = 16'h3cc7; 14'h a8b: x = 16'h3cc6; 14'h a8c: x = 16'h3cc4; 14'h a8d: x = 16'h3cc2; 14'h a8e: x = 16'h3cc1; 14'h a8f: x = 16'h3cbf; 14'h a90: x = 16'h3cbe; 14'h a91: x = 16'h3cbc; 14'h a92: x = 16'h3cba; 14'h a93: x = 16'h3cb9; 14'h a94: x = 16'h3cb7; 14'h a95: x = 16'h3cb6; 14'h a96: x = 16'h3cb4; 14'h a97: x = 16'h3cb2; 14'h a98: x = 16'h3cb1; 14'h a99: x = 16'h3caf; 14'h a9a: x = 16'h3cae; 14'h a9b: x = 16'h3cac; 14'h a9c: x = 16'h3caa; 14'h a9d: x = 16'h3ca9; 14'h a9e: x = 16'h3ca7; 14'h a9f: x = 16'h3ca6; 14'h aa0: x = 16'h3ca4; 14'h aa1: x = 16'h3ca2; 14'h aa2: x = 16'h3ca1; 14'h aa3: x = 16'h3c9f; 14'h aa4: x = 16'h3c9e; 14'h aa5: x = 16'h3c9c; 14'h aa6: x = 16'h3c9b; 14'h aa7: x = 16'h3c99; 14'h aa8: x = 16'h3c97; 14'h aa9: x = 16'h3c96; 14'h aaa: x = 16'h3c94; 14'h aab: x = 16'h3c93; 14'h aac: x = 16'h3c91; 14'h aad: x = 16'h3c8f; 14'h aae: x = 16'h3c8e; 14'h aaf: x = 16'h3c8c; 14'h ab0: x = 16'h3c8b; 14'h ab1: x = 16'h3c89; 14'h ab2: x = 16'h3c87; 14'h ab3: x = 16'h3c86; 14'h ab4: x = 16'h3c84; 14'h ab5: x = 16'h3c83; 14'h ab6: x = 16'h3c81; 14'h ab7: x = 16'h3c80; 14'h ab8: x = 16'h3c7e; 14'h ab9: x = 16'h3c7c; 14'h aba: x = 16'h3c7b; 14'h abb: x = 16'h3c79; 14'h abc: x = 16'h3c78; 14'h abd: x = 16'h3c76; 14'h abe: x = 16'h3c75; 14'h abf: x = 16'h3c73; 14'h ac0: x = 16'h3c71; 14'h ac1: x = 16'h3c70; 14'h ac2: x = 16'h3c6e; 14'h ac3: x = 16'h3c6d; 14'h ac4: x = 16'h3c6b; 14'h ac5: x = 16'h3c6a; 14'h ac6: x = 16'h3c68; 14'h ac7: x = 16'h3c66; 14'h ac8: x = 16'h3c65; 14'h ac9: x = 16'h3c63; 14'h aca: x = 16'h3c62; 14'h acb: x = 16'h3c60; 14'h acc: x = 16'h3c5f; 14'h acd: x = 16'h3c5d; 14'h ace: x = 16'h3c5b; 14'h acf: x = 16'h3c5a; 14'h ad0: x = 16'h3c58; 14'h ad1: x = 16'h3c57; 14'h ad2: x = 16'h3c55; 14'h ad3: x = 16'h3c54; 14'h ad4: x = 16'h3c52; 14'h ad5: x = 16'h3c50; 14'h ad6: x = 16'h3c4f; 14'h ad7: x = 16'h3c4d; 14'h ad8: x = 16'h3c4c; 14'h ad9: x = 16'h3c4a; 14'h ada: x = 16'h3c49; 14'h adb: x = 16'h3c47; 14'h adc: x = 16'h3c45; 14'h add: x = 16'h3c44; 14'h ade: x = 16'h3c42; 14'h adf: x = 16'h3c41; 14'h ae0: x = 16'h3c3f; 14'h ae1: x = 16'h3c3e; 14'h ae2: x = 16'h3c3c; 14'h ae3: x = 16'h3c3a; 14'h ae4: x = 16'h3c39; 14'h ae5: x = 16'h3c37; 14'h ae6: x = 16'h3c36; 14'h ae7: x = 16'h3c34; 14'h ae8: x = 16'h3c33; 14'h ae9: x = 16'h3c31; 14'h aea: x = 16'h3c30; 14'h aeb: x = 16'h3c2e; 14'h aec: x = 16'h3c2c; 14'h aed: x = 16'h3c2b; 14'h aee: x = 16'h3c29; 14'h aef: x = 16'h3c28; 14'h af0: x = 16'h3c26; 14'h af1: x = 16'h3c25; 14'h af2: x = 16'h3c23; 14'h af3: x = 16'h3c22; 14'h af4: x = 16'h3c20; 14'h af5: x = 16'h3c1e; 14'h af6: x = 16'h3c1d; 14'h af7: x = 16'h3c1b; 14'h af8: x = 16'h3c1a; 14'h af9: x = 16'h3c18; 14'h afa: x = 16'h3c17; 14'h afb: x = 16'h3c15; 14'h afc: x = 16'h3c14; 14'h afd: x = 16'h3c12; 14'h afe: x = 16'h3c10; 14'h aff: x = 16'h3c0f; 14'h b00: x = 16'h3c0d; 14'h b01: x = 16'h3c0c; 14'h b02: x = 16'h3c0a; 14'h b03: x = 16'h3c09; 14'h b04: x = 16'h3c07; 14'h b05: x = 16'h3c06; 14'h b06: x = 16'h3c04; 14'h b07: x = 16'h3c03; 14'h b08: x = 16'h3c01; 14'h b09: x = 16'h3bff; 14'h b0a: x = 16'h3bfe; 14'h b0b: x = 16'h3bfc; 14'h b0c: x = 16'h3bfb; 14'h b0d: x = 16'h3bf9; 14'h b0e: x = 16'h3bf8; 14'h b0f: x = 16'h3bf6; 14'h b10: x = 16'h3bf5; 14'h b11: x = 16'h3bf3; 14'h b12: x = 16'h3bf2; 14'h b13: x = 16'h3bf0; 14'h b14: x = 16'h3bee; 14'h b15: x = 16'h3bed; 14'h b16: x = 16'h3beb; 14'h b17: x = 16'h3bea; 14'h b18: x = 16'h3be8; 14'h b19: x = 16'h3be7; 14'h b1a: x = 16'h3be5; 14'h b1b: x = 16'h3be4; 14'h b1c: x = 16'h3be2; 14'h b1d: x = 16'h3be1; 14'h b1e: x = 16'h3bdf; 14'h b1f: x = 16'h3bde; 14'h b20: x = 16'h3bdc; 14'h b21: x = 16'h3bda; 14'h b22: x = 16'h3bd9; 14'h b23: x = 16'h3bd7; 14'h b24: x = 16'h3bd6; 14'h b25: x = 16'h3bd4; 14'h b26: x = 16'h3bd3; 14'h b27: x = 16'h3bd1; 14'h b28: x = 16'h3bd0; 14'h b29: x = 16'h3bce; 14'h b2a: x = 16'h3bcd; 14'h b2b: x = 16'h3bcb; 14'h b2c: x = 16'h3bca; 14'h b2d: x = 16'h3bc8; 14'h b2e: x = 16'h3bc6; 14'h b2f: x = 16'h3bc5; 14'h b30: x = 16'h3bc3; 14'h b31: x = 16'h3bc2; 14'h b32: x = 16'h3bc0; 14'h b33: x = 16'h3bbf; 14'h b34: x = 16'h3bbd; 14'h b35: x = 16'h3bbc; 14'h b36: x = 16'h3bba; 14'h b37: x = 16'h3bb9; 14'h b38: x = 16'h3bb7; 14'h b39: x = 16'h3bb6; 14'h b3a: x = 16'h3bb4; 14'h b3b: x = 16'h3bb3; 14'h b3c: x = 16'h3bb1; 14'h b3d: x = 16'h3bb0; 14'h b3e: x = 16'h3bae; 14'h b3f: x = 16'h3bac; 14'h b40: x = 16'h3bab; 14'h b41: x = 16'h3ba9; 14'h b42: x = 16'h3ba8; 14'h b43: x = 16'h3ba6; 14'h b44: x = 16'h3ba5; 14'h b45: x = 16'h3ba3; 14'h b46: x = 16'h3ba2; 14'h b47: x = 16'h3ba0; 14'h b48: x = 16'h3b9f; 14'h b49: x = 16'h3b9d; 14'h b4a: x = 16'h3b9c; 14'h b4b: x = 16'h3b9a; 14'h b4c: x = 16'h3b99; 14'h b4d: x = 16'h3b97; 14'h b4e: x = 16'h3b96; 14'h b4f: x = 16'h3b94; 14'h b50: x = 16'h3b93; 14'h b51: x = 16'h3b91; 14'h b52: x = 16'h3b90; 14'h b53: x = 16'h3b8e; 14'h b54: x = 16'h3b8d; 14'h b55: x = 16'h3b8b; 14'h b56: x = 16'h3b89; 14'h b57: x = 16'h3b88; 14'h b58: x = 16'h3b86; 14'h b59: x = 16'h3b85; 14'h b5a: x = 16'h3b83; 14'h b5b: x = 16'h3b82; 14'h b5c: x = 16'h3b80; 14'h b5d: x = 16'h3b7f; 14'h b5e: x = 16'h3b7d; 14'h b5f: x = 16'h3b7c; 14'h b60: x = 16'h3b7a; 14'h b61: x = 16'h3b79; 14'h b62: x = 16'h3b77; 14'h b63: x = 16'h3b76; 14'h b64: x = 16'h3b74; 14'h b65: x = 16'h3b73; 14'h b66: x = 16'h3b71; 14'h b67: x = 16'h3b70; 14'h b68: x = 16'h3b6e; 14'h b69: x = 16'h3b6d; 14'h b6a: x = 16'h3b6b; 14'h b6b: x = 16'h3b6a; 14'h b6c: x = 16'h3b68; 14'h b6d: x = 16'h3b67; 14'h b6e: x = 16'h3b65; 14'h b6f: x = 16'h3b64; 14'h b70: x = 16'h3b62; 14'h b71: x = 16'h3b61; 14'h b72: x = 16'h3b5f; 14'h b73: x = 16'h3b5e; 14'h b74: x = 16'h3b5c; 14'h b75: x = 16'h3b5b; 14'h b76: x = 16'h3b59; 14'h b77: x = 16'h3b58; 14'h b78: x = 16'h3b56; 14'h b79: x = 16'h3b55; 14'h b7a: x = 16'h3b53; 14'h b7b: x = 16'h3b52; 14'h b7c: x = 16'h3b50; 14'h b7d: x = 16'h3b4f; 14'h b7e: x = 16'h3b4d; 14'h b7f: x = 16'h3b4c; 14'h b80: x = 16'h3b4a; 14'h b81: x = 16'h3b49; 14'h b82: x = 16'h3b47; 14'h b83: x = 16'h3b46; 14'h b84: x = 16'h3b44; 14'h b85: x = 16'h3b43; 14'h b86: x = 16'h3b41; 14'h b87: x = 16'h3b40; 14'h b88: x = 16'h3b3e; 14'h b89: x = 16'h3b3d; 14'h b8a: x = 16'h3b3b; 14'h b8b: x = 16'h3b3a; 14'h b8c: x = 16'h3b38; 14'h b8d: x = 16'h3b37; 14'h b8e: x = 16'h3b35; 14'h b8f: x = 16'h3b34; 14'h b90: x = 16'h3b32; 14'h b91: x = 16'h3b31; 14'h b92: x = 16'h3b2f; 14'h b93: x = 16'h3b2e; 14'h b94: x = 16'h3b2c; 14'h b95: x = 16'h3b2b; 14'h b96: x = 16'h3b29; 14'h b97: x = 16'h3b28; 14'h b98: x = 16'h3b26; 14'h b99: x = 16'h3b25; 14'h b9a: x = 16'h3b23; 14'h b9b: x = 16'h3b22; 14'h b9c: x = 16'h3b20; 14'h b9d: x = 16'h3b1f; 14'h b9e: x = 16'h3b1d; 14'h b9f: x = 16'h3b1c; 14'h ba0: x = 16'h3b1a; 14'h ba1: x = 16'h3b19; 14'h ba2: x = 16'h3b17; 14'h ba3: x = 16'h3b16; 14'h ba4: x = 16'h3b14; 14'h ba5: x = 16'h3b13; 14'h ba6: x = 16'h3b11; 14'h ba7: x = 16'h3b10; 14'h ba8: x = 16'h3b0e; 14'h ba9: x = 16'h3b0d; 14'h baa: x = 16'h3b0b; 14'h bab: x = 16'h3b0a; 14'h bac: x = 16'h3b08; 14'h bad: x = 16'h3b07; 14'h bae: x = 16'h3b05; 14'h baf: x = 16'h3b04; 14'h bb0: x = 16'h3b02; 14'h bb1: x = 16'h3b01; 14'h bb2: x = 16'h3aff; 14'h bb3: x = 16'h3afe; 14'h bb4: x = 16'h3afc; 14'h bb5: x = 16'h3afb; 14'h bb6: x = 16'h3afa; 14'h bb7: x = 16'h3af8; 14'h bb8: x = 16'h3af7; 14'h bb9: x = 16'h3af5; 14'h bba: x = 16'h3af4; 14'h bbb: x = 16'h3af2; 14'h bbc: x = 16'h3af1; 14'h bbd: x = 16'h3aef; 14'h bbe: x = 16'h3aee; 14'h bbf: x = 16'h3aec; 14'h bc0: x = 16'h3aeb; 14'h bc1: x = 16'h3ae9; 14'h bc2: x = 16'h3ae8; 14'h bc3: x = 16'h3ae6; 14'h bc4: x = 16'h3ae5; 14'h bc5: x = 16'h3ae3; 14'h bc6: x = 16'h3ae2; 14'h bc7: x = 16'h3ae0; 14'h bc8: x = 16'h3adf; 14'h bc9: x = 16'h3add; 14'h bca: x = 16'h3adc; 14'h bcb: x = 16'h3ada; 14'h bcc: x = 16'h3ad9; 14'h bcd: x = 16'h3ad8; 14'h bce: x = 16'h3ad6; 14'h bcf: x = 16'h3ad5; 14'h bd0: x = 16'h3ad3; 14'h bd1: x = 16'h3ad2; 14'h bd2: x = 16'h3ad0; 14'h bd3: x = 16'h3acf; 14'h bd4: x = 16'h3acd; 14'h bd5: x = 16'h3acc; 14'h bd6: x = 16'h3aca; 14'h bd7: x = 16'h3ac9; 14'h bd8: x = 16'h3ac7; 14'h bd9: x = 16'h3ac6; 14'h bda: x = 16'h3ac4; 14'h bdb: x = 16'h3ac3; 14'h bdc: x = 16'h3ac1; 14'h bdd: x = 16'h3ac0; 14'h bde: x = 16'h3abe; 14'h bdf: x = 16'h3abd; 14'h be0: x = 16'h3abc; 14'h be1: x = 16'h3aba; 14'h be2: x = 16'h3ab9; 14'h be3: x = 16'h3ab7; 14'h be4: x = 16'h3ab6; 14'h be5: x = 16'h3ab4; 14'h be6: x = 16'h3ab3; 14'h be7: x = 16'h3ab1; 14'h be8: x = 16'h3ab0; 14'h be9: x = 16'h3aae; 14'h bea: x = 16'h3aad; 14'h beb: x = 16'h3aab; 14'h bec: x = 16'h3aaa; 14'h bed: x = 16'h3aa8; 14'h bee: x = 16'h3aa7; 14'h bef: x = 16'h3aa6; 14'h bf0: x = 16'h3aa4; 14'h bf1: x = 16'h3aa3; 14'h bf2: x = 16'h3aa1; 14'h bf3: x = 16'h3aa0; 14'h bf4: x = 16'h3a9e; 14'h bf5: x = 16'h3a9d; 14'h bf6: x = 16'h3a9b; 14'h bf7: x = 16'h3a9a; 14'h bf8: x = 16'h3a98; 14'h bf9: x = 16'h3a97; 14'h bfa: x = 16'h3a95; 14'h bfb: x = 16'h3a94; 14'h bfc: x = 16'h3a93; 14'h bfd: x = 16'h3a91; 14'h bfe: x = 16'h3a90; 14'h bff: x = 16'h3a8e; 14'h c00: x = 16'h3a8d; 14'h c01: x = 16'h3a8b; 14'h c02: x = 16'h3a8a; 14'h c03: x = 16'h3a88; 14'h c04: x = 16'h3a87; 14'h c05: x = 16'h3a85; 14'h c06: x = 16'h3a84; 14'h c07: x = 16'h3a83; 14'h c08: x = 16'h3a81; 14'h c09: x = 16'h3a80; 14'h c0a: x = 16'h3a7e; 14'h c0b: x = 16'h3a7d; 14'h c0c: x = 16'h3a7b; 14'h c0d: x = 16'h3a7a; 14'h c0e: x = 16'h3a78; 14'h c0f: x = 16'h3a77; 14'h c10: x = 16'h3a75; 14'h c11: x = 16'h3a74; 14'h c12: x = 16'h3a73; 14'h c13: x = 16'h3a71; 14'h c14: x = 16'h3a70; 14'h c15: x = 16'h3a6e; 14'h c16: x = 16'h3a6d; 14'h c17: x = 16'h3a6b; 14'h c18: x = 16'h3a6a; 14'h c19: x = 16'h3a68; 14'h c1a: x = 16'h3a67; 14'h c1b: x = 16'h3a66; 14'h c1c: x = 16'h3a64; 14'h c1d: x = 16'h3a63; 14'h c1e: x = 16'h3a61; 14'h c1f: x = 16'h3a60; 14'h c20: x = 16'h3a5e; 14'h c21: x = 16'h3a5d; 14'h c22: x = 16'h3a5b; 14'h c23: x = 16'h3a5a; 14'h c24: x = 16'h3a58; 14'h c25: x = 16'h3a57; 14'h c26: x = 16'h3a56; 14'h c27: x = 16'h3a54; 14'h c28: x = 16'h3a53; 14'h c29: x = 16'h3a51; 14'h c2a: x = 16'h3a50; 14'h c2b: x = 16'h3a4e; 14'h c2c: x = 16'h3a4d; 14'h c2d: x = 16'h3a4b; 14'h c2e: x = 16'h3a4a; 14'h c2f: x = 16'h3a49; 14'h c30: x = 16'h3a47; 14'h c31: x = 16'h3a46; 14'h c32: x = 16'h3a44; 14'h c33: x = 16'h3a43; 14'h c34: x = 16'h3a41; 14'h c35: x = 16'h3a40; 14'h c36: x = 16'h3a3f; 14'h c37: x = 16'h3a3d; 14'h c38: x = 16'h3a3c; 14'h c39: x = 16'h3a3a; 14'h c3a: x = 16'h3a39; 14'h c3b: x = 16'h3a37; 14'h c3c: x = 16'h3a36; 14'h c3d: x = 16'h3a34; 14'h c3e: x = 16'h3a33; 14'h c3f: x = 16'h3a32; 14'h c40: x = 16'h3a30; 14'h c41: x = 16'h3a2f; 14'h c42: x = 16'h3a2d; 14'h c43: x = 16'h3a2c; 14'h c44: x = 16'h3a2a; 14'h c45: x = 16'h3a29; 14'h c46: x = 16'h3a28; 14'h c47: x = 16'h3a26; 14'h c48: x = 16'h3a25; 14'h c49: x = 16'h3a23; 14'h c4a: x = 16'h3a22; 14'h c4b: x = 16'h3a20; 14'h c4c: x = 16'h3a1f; 14'h c4d: x = 16'h3a1d; 14'h c4e: x = 16'h3a1c; 14'h c4f: x = 16'h3a1b; 14'h c50: x = 16'h3a19; 14'h c51: x = 16'h3a18; 14'h c52: x = 16'h3a16; 14'h c53: x = 16'h3a15; 14'h c54: x = 16'h3a13; 14'h c55: x = 16'h3a12; 14'h c56: x = 16'h3a11; 14'h c57: x = 16'h3a0f; 14'h c58: x = 16'h3a0e; 14'h c59: x = 16'h3a0c; 14'h c5a: x = 16'h3a0b; 14'h c5b: x = 16'h3a09; 14'h c5c: x = 16'h3a08; 14'h c5d: x = 16'h3a07; 14'h c5e: x = 16'h3a05; 14'h c5f: x = 16'h3a04; 14'h c60: x = 16'h3a02; 14'h c61: x = 16'h3a01; 14'h c62: x = 16'h39ff; 14'h c63: x = 16'h39fe; 14'h c64: x = 16'h39fd; 14'h c65: x = 16'h39fb; 14'h c66: x = 16'h39fa; 14'h c67: x = 16'h39f8; 14'h c68: x = 16'h39f7; 14'h c69: x = 16'h39f6; 14'h c6a: x = 16'h39f4; 14'h c6b: x = 16'h39f3; 14'h c6c: x = 16'h39f1; 14'h c6d: x = 16'h39f0; 14'h c6e: x = 16'h39ee; 14'h c6f: x = 16'h39ed; 14'h c70: x = 16'h39ec; 14'h c71: x = 16'h39ea; 14'h c72: x = 16'h39e9; 14'h c73: x = 16'h39e7; 14'h c74: x = 16'h39e6; 14'h c75: x = 16'h39e4; 14'h c76: x = 16'h39e3; 14'h c77: x = 16'h39e2; 14'h c78: x = 16'h39e0; 14'h c79: x = 16'h39df; 14'h c7a: x = 16'h39dd; 14'h c7b: x = 16'h39dc; 14'h c7c: x = 16'h39db; 14'h c7d: x = 16'h39d9; 14'h c7e: x = 16'h39d8; 14'h c7f: x = 16'h39d6; 14'h c80: x = 16'h39d5; 14'h c81: x = 16'h39d3; 14'h c82: x = 16'h39d2; 14'h c83: x = 16'h39d1; 14'h c84: x = 16'h39cf; 14'h c85: x = 16'h39ce; 14'h c86: x = 16'h39cc; 14'h c87: x = 16'h39cb; 14'h c88: x = 16'h39ca; 14'h c89: x = 16'h39c8; 14'h c8a: x = 16'h39c7; 14'h c8b: x = 16'h39c5; 14'h c8c: x = 16'h39c4; 14'h c8d: x = 16'h39c2; 14'h c8e: x = 16'h39c1; 14'h c8f: x = 16'h39c0; 14'h c90: x = 16'h39be; 14'h c91: x = 16'h39bd; 14'h c92: x = 16'h39bb; 14'h c93: x = 16'h39ba; 14'h c94: x = 16'h39b9; 14'h c95: x = 16'h39b7; 14'h c96: x = 16'h39b6; 14'h c97: x = 16'h39b4; 14'h c98: x = 16'h39b3; 14'h c99: x = 16'h39b2; 14'h c9a: x = 16'h39b0; 14'h c9b: x = 16'h39af; 14'h c9c: x = 16'h39ad; 14'h c9d: x = 16'h39ac; 14'h c9e: x = 16'h39aa; 14'h c9f: x = 16'h39a9; 14'h ca0: x = 16'h39a8; 14'h ca1: x = 16'h39a6; 14'h ca2: x = 16'h39a5; 14'h ca3: x = 16'h39a3; 14'h ca4: x = 16'h39a2; 14'h ca5: x = 16'h39a1; 14'h ca6: x = 16'h399f; 14'h ca7: x = 16'h399e; 14'h ca8: x = 16'h399c; 14'h ca9: x = 16'h399b; 14'h caa: x = 16'h399a; 14'h cab: x = 16'h3998; 14'h cac: x = 16'h3997; 14'h cad: x = 16'h3995; 14'h cae: x = 16'h3994; 14'h caf: x = 16'h3993; 14'h cb0: x = 16'h3991; 14'h cb1: x = 16'h3990; 14'h cb2: x = 16'h398e; 14'h cb3: x = 16'h398d; 14'h cb4: x = 16'h398c; 14'h cb5: x = 16'h398a; 14'h cb6: x = 16'h3989; 14'h cb7: x = 16'h3987; 14'h cb8: x = 16'h3986; 14'h cb9: x = 16'h3985; 14'h cba: x = 16'h3983; 14'h cbb: x = 16'h3982; 14'h cbc: x = 16'h3980; 14'h cbd: x = 16'h397f; 14'h cbe: x = 16'h397e; 14'h cbf: x = 16'h397c; 14'h cc0: x = 16'h397b; 14'h cc1: x = 16'h3979; 14'h cc2: x = 16'h3978; 14'h cc3: x = 16'h3977; 14'h cc4: x = 16'h3975; 14'h cc5: x = 16'h3974; 14'h cc6: x = 16'h3972; 14'h cc7: x = 16'h3971; 14'h cc8: x = 16'h3970; 14'h cc9: x = 16'h396e; 14'h cca: x = 16'h396d; 14'h ccb: x = 16'h396b; 14'h ccc: x = 16'h396a; 14'h ccd: x = 16'h3969; 14'h cce: x = 16'h3967; 14'h ccf: x = 16'h3966; 14'h cd0: x = 16'h3964; 14'h cd1: x = 16'h3963; 14'h cd2: x = 16'h3962; 14'h cd3: x = 16'h3960; 14'h cd4: x = 16'h395f; 14'h cd5: x = 16'h395e; 14'h cd6: x = 16'h395c; 14'h cd7: x = 16'h395b; 14'h cd8: x = 16'h3959; 14'h cd9: x = 16'h3958; 14'h cda: x = 16'h3957; 14'h cdb: x = 16'h3955; 14'h cdc: x = 16'h3954; 14'h cdd: x = 16'h3952; 14'h cde: x = 16'h3951; 14'h cdf: x = 16'h3950; 14'h ce0: x = 16'h394e; 14'h ce1: x = 16'h394d; 14'h ce2: x = 16'h394b; 14'h ce3: x = 16'h394a; 14'h ce4: x = 16'h3949; 14'h ce5: x = 16'h3947; 14'h ce6: x = 16'h3946; 14'h ce7: x = 16'h3945; 14'h ce8: x = 16'h3943; 14'h ce9: x = 16'h3942; 14'h cea: x = 16'h3940; 14'h ceb: x = 16'h393f; 14'h cec: x = 16'h393e; 14'h ced: x = 16'h393c; 14'h cee: x = 16'h393b; 14'h cef: x = 16'h3939; 14'h cf0: x = 16'h3938; 14'h cf1: x = 16'h3937; 14'h cf2: x = 16'h3935; 14'h cf3: x = 16'h3934; 14'h cf4: x = 16'h3933; 14'h cf5: x = 16'h3931; 14'h cf6: x = 16'h3930; 14'h cf7: x = 16'h392e; 14'h cf8: x = 16'h392d; 14'h cf9: x = 16'h392c; 14'h cfa: x = 16'h392a; 14'h cfb: x = 16'h3929; 14'h cfc: x = 16'h3928; 14'h cfd: x = 16'h3926; 14'h cfe: x = 16'h3925; 14'h cff: x = 16'h3923; 14'h d00: x = 16'h3922; 14'h d01: x = 16'h3921; 14'h d02: x = 16'h391f; 14'h d03: x = 16'h391e; 14'h d04: x = 16'h391c; 14'h d05: x = 16'h391b; 14'h d06: x = 16'h391a; 14'h d07: x = 16'h3918; 14'h d08: x = 16'h3917; 14'h d09: x = 16'h3916; 14'h d0a: x = 16'h3914; 14'h d0b: x = 16'h3913; 14'h d0c: x = 16'h3911; 14'h d0d: x = 16'h3910; 14'h d0e: x = 16'h390f; 14'h d0f: x = 16'h390d; 14'h d10: x = 16'h390c; 14'h d11: x = 16'h390b; 14'h d12: x = 16'h3909; 14'h d13: x = 16'h3908; 14'h d14: x = 16'h3906; 14'h d15: x = 16'h3905; 14'h d16: x = 16'h3904; 14'h d17: x = 16'h3902; 14'h d18: x = 16'h3901; 14'h d19: x = 16'h3900; 14'h d1a: x = 16'h38fe; 14'h d1b: x = 16'h38fd; 14'h d1c: x = 16'h38fb; 14'h d1d: x = 16'h38fa; 14'h d1e: x = 16'h38f9; 14'h d1f: x = 16'h38f7; 14'h d20: x = 16'h38f6; 14'h d21: x = 16'h38f5; 14'h d22: x = 16'h38f3; 14'h d23: x = 16'h38f2; 14'h d24: x = 16'h38f1; 14'h d25: x = 16'h38ef; 14'h d26: x = 16'h38ee; 14'h d27: x = 16'h38ec; 14'h d28: x = 16'h38eb; 14'h d29: x = 16'h38ea; 14'h d2a: x = 16'h38e8; 14'h d2b: x = 16'h38e7; 14'h d2c: x = 16'h38e6; 14'h d2d: x = 16'h38e4; 14'h d2e: x = 16'h38e3; 14'h d2f: x = 16'h38e2; 14'h d30: x = 16'h38e0; 14'h d31: x = 16'h38df; 14'h d32: x = 16'h38dd; 14'h d33: x = 16'h38dc; 14'h d34: x = 16'h38db; 14'h d35: x = 16'h38d9; 14'h d36: x = 16'h38d8; 14'h d37: x = 16'h38d7; 14'h d38: x = 16'h38d5; 14'h d39: x = 16'h38d4; 14'h d3a: x = 16'h38d2; 14'h d3b: x = 16'h38d1; 14'h d3c: x = 16'h38d0; 14'h d3d: x = 16'h38ce; 14'h d3e: x = 16'h38cd; 14'h d3f: x = 16'h38cc; 14'h d40: x = 16'h38ca; 14'h d41: x = 16'h38c9; 14'h d42: x = 16'h38c8; 14'h d43: x = 16'h38c6; 14'h d44: x = 16'h38c5; 14'h d45: x = 16'h38c4; 14'h d46: x = 16'h38c2; 14'h d47: x = 16'h38c1; 14'h d48: x = 16'h38bf; 14'h d49: x = 16'h38be; 14'h d4a: x = 16'h38bd; 14'h d4b: x = 16'h38bb; 14'h d4c: x = 16'h38ba; 14'h d4d: x = 16'h38b9; 14'h d4e: x = 16'h38b7; 14'h d4f: x = 16'h38b6; 14'h d50: x = 16'h38b5; 14'h d51: x = 16'h38b3; 14'h d52: x = 16'h38b2; 14'h d53: x = 16'h38b1; 14'h d54: x = 16'h38af; 14'h d55: x = 16'h38ae; 14'h d56: x = 16'h38ac; 14'h d57: x = 16'h38ab; 14'h d58: x = 16'h38aa; 14'h d59: x = 16'h38a8; 14'h d5a: x = 16'h38a7; 14'h d5b: x = 16'h38a6; 14'h d5c: x = 16'h38a4; 14'h d5d: x = 16'h38a3; 14'h d5e: x = 16'h38a2; 14'h d5f: x = 16'h38a0; 14'h d60: x = 16'h389f; 14'h d61: x = 16'h389e; 14'h d62: x = 16'h389c; 14'h d63: x = 16'h389b; 14'h d64: x = 16'h389a; 14'h d65: x = 16'h3898; 14'h d66: x = 16'h3897; 14'h d67: x = 16'h3895; 14'h d68: x = 16'h3894; 14'h d69: x = 16'h3893; 14'h d6a: x = 16'h3891; 14'h d6b: x = 16'h3890; 14'h d6c: x = 16'h388f; 14'h d6d: x = 16'h388d; 14'h d6e: x = 16'h388c; 14'h d6f: x = 16'h388b; 14'h d70: x = 16'h3889; 14'h d71: x = 16'h3888; 14'h d72: x = 16'h3887; 14'h d73: x = 16'h3885; 14'h d74: x = 16'h3884; 14'h d75: x = 16'h3883; 14'h d76: x = 16'h3881; 14'h d77: x = 16'h3880; 14'h d78: x = 16'h387f; 14'h d79: x = 16'h387d; 14'h d7a: x = 16'h387c; 14'h d7b: x = 16'h387b; 14'h d7c: x = 16'h3879; 14'h d7d: x = 16'h3878; 14'h d7e: x = 16'h3876; 14'h d7f: x = 16'h3875; 14'h d80: x = 16'h3874; 14'h d81: x = 16'h3872; 14'h d82: x = 16'h3871; 14'h d83: x = 16'h3870; 14'h d84: x = 16'h386e; 14'h d85: x = 16'h386d; 14'h d86: x = 16'h386c; 14'h d87: x = 16'h386a; 14'h d88: x = 16'h3869; 14'h d89: x = 16'h3868; 14'h d8a: x = 16'h3866; 14'h d8b: x = 16'h3865; 14'h d8c: x = 16'h3864; 14'h d8d: x = 16'h3862; 14'h d8e: x = 16'h3861; 14'h d8f: x = 16'h3860; 14'h d90: x = 16'h385e; 14'h d91: x = 16'h385d; 14'h d92: x = 16'h385c; 14'h d93: x = 16'h385a; 14'h d94: x = 16'h3859; 14'h d95: x = 16'h3858; 14'h d96: x = 16'h3856; 14'h d97: x = 16'h3855; 14'h d98: x = 16'h3854; 14'h d99: x = 16'h3852; 14'h d9a: x = 16'h3851; 14'h d9b: x = 16'h3850; 14'h d9c: x = 16'h384e; 14'h d9d: x = 16'h384d; 14'h d9e: x = 16'h384c; 14'h d9f: x = 16'h384a; 14'h da0: x = 16'h3849; 14'h da1: x = 16'h3848; 14'h da2: x = 16'h3846; 14'h da3: x = 16'h3845; 14'h da4: x = 16'h3844; 14'h da5: x = 16'h3842; 14'h da6: x = 16'h3841; 14'h da7: x = 16'h3840; 14'h da8: x = 16'h383e; 14'h da9: x = 16'h383d; 14'h daa: x = 16'h383c; 14'h dab: x = 16'h383a; 14'h dac: x = 16'h3839; 14'h dad: x = 16'h3838; 14'h dae: x = 16'h3836; 14'h daf: x = 16'h3835; 14'h db0: x = 16'h3834; 14'h db1: x = 16'h3832; 14'h db2: x = 16'h3831; 14'h db3: x = 16'h3830; 14'h db4: x = 16'h382e; 14'h db5: x = 16'h382d; 14'h db6: x = 16'h382c; 14'h db7: x = 16'h382a; 14'h db8: x = 16'h3829; 14'h db9: x = 16'h3828; 14'h dba: x = 16'h3826; 14'h dbb: x = 16'h3825; 14'h dbc: x = 16'h3824; 14'h dbd: x = 16'h3822; 14'h dbe: x = 16'h3821; 14'h dbf: x = 16'h3820; 14'h dc0: x = 16'h381e; 14'h dc1: x = 16'h381d; 14'h dc2: x = 16'h381c; 14'h dc3: x = 16'h381a; 14'h dc4: x = 16'h3819; 14'h dc5: x = 16'h3818; 14'h dc6: x = 16'h3816; 14'h dc7: x = 16'h3815; 14'h dc8: x = 16'h3814; 14'h dc9: x = 16'h3812; 14'h dca: x = 16'h3811; 14'h dcb: x = 16'h3810; 14'h dcc: x = 16'h380e; 14'h dcd: x = 16'h380d; 14'h dce: x = 16'h380c; 14'h dcf: x = 16'h380a; 14'h dd0: x = 16'h3809; 14'h dd1: x = 16'h3808; 14'h dd2: x = 16'h3806; 14'h dd3: x = 16'h3805; 14'h dd4: x = 16'h3804; 14'h dd5: x = 16'h3803; 14'h dd6: x = 16'h3801; 14'h dd7: x = 16'h3800; 14'h dd8: x = 16'h37ff; 14'h dd9: x = 16'h37fd; 14'h dda: x = 16'h37fc; 14'h ddb: x = 16'h37fb; 14'h ddc: x = 16'h37f9; 14'h ddd: x = 16'h37f8; 14'h dde: x = 16'h37f7; 14'h ddf: x = 16'h37f5; 14'h de0: x = 16'h37f4; 14'h de1: x = 16'h37f3; 14'h de2: x = 16'h37f1; 14'h de3: x = 16'h37f0; 14'h de4: x = 16'h37ef; 14'h de5: x = 16'h37ed; 14'h de6: x = 16'h37ec; 14'h de7: x = 16'h37eb; 14'h de8: x = 16'h37e9; 14'h de9: x = 16'h37e8; 14'h dea: x = 16'h37e7; 14'h deb: x = 16'h37e6; 14'h dec: x = 16'h37e4; 14'h ded: x = 16'h37e3; 14'h dee: x = 16'h37e2; 14'h def: x = 16'h37e0; 14'h df0: x = 16'h37df; 14'h df1: x = 16'h37de; 14'h df2: x = 16'h37dc; 14'h df3: x = 16'h37db; 14'h df4: x = 16'h37da; 14'h df5: x = 16'h37d8; 14'h df6: x = 16'h37d7; 14'h df7: x = 16'h37d6; 14'h df8: x = 16'h37d4; 14'h df9: x = 16'h37d3; 14'h dfa: x = 16'h37d2; 14'h dfb: x = 16'h37d0; 14'h dfc: x = 16'h37cf; 14'h dfd: x = 16'h37ce; 14'h dfe: x = 16'h37cd; 14'h dff: x = 16'h37cb; 14'h e00: x = 16'h37ca; 14'h e01: x = 16'h37c9; 14'h e02: x = 16'h37c7; 14'h e03: x = 16'h37c6; 14'h e04: x = 16'h37c5; 14'h e05: x = 16'h37c3; 14'h e06: x = 16'h37c2; 14'h e07: x = 16'h37c1; 14'h e08: x = 16'h37bf; 14'h e09: x = 16'h37be; 14'h e0a: x = 16'h37bd; 14'h e0b: x = 16'h37bc; 14'h e0c: x = 16'h37ba; 14'h e0d: x = 16'h37b9; 14'h e0e: x = 16'h37b8; 14'h e0f: x = 16'h37b6; 14'h e10: x = 16'h37b5; 14'h e11: x = 16'h37b4; 14'h e12: x = 16'h37b2; 14'h e13: x = 16'h37b1; 14'h e14: x = 16'h37b0; 14'h e15: x = 16'h37ae; 14'h e16: x = 16'h37ad; 14'h e17: x = 16'h37ac; 14'h e18: x = 16'h37ab; 14'h e19: x = 16'h37a9; 14'h e1a: x = 16'h37a8; 14'h e1b: x = 16'h37a7; 14'h e1c: x = 16'h37a5; 14'h e1d: x = 16'h37a4; 14'h e1e: x = 16'h37a3; 14'h e1f: x = 16'h37a1; 14'h e20: x = 16'h37a0; 14'h e21: x = 16'h379f; 14'h e22: x = 16'h379d; 14'h e23: x = 16'h379c; 14'h e24: x = 16'h379b; 14'h e25: x = 16'h379a; 14'h e26: x = 16'h3798; 14'h e27: x = 16'h3797; 14'h e28: x = 16'h3796; 14'h e29: x = 16'h3794; 14'h e2a: x = 16'h3793; 14'h e2b: x = 16'h3792; 14'h e2c: x = 16'h3790; 14'h e2d: x = 16'h378f; 14'h e2e: x = 16'h378e; 14'h e2f: x = 16'h378d; 14'h e30: x = 16'h378b; 14'h e31: x = 16'h378a; 14'h e32: x = 16'h3789; 14'h e33: x = 16'h3787; 14'h e34: x = 16'h3786; 14'h e35: x = 16'h3785; 14'h e36: x = 16'h3783; 14'h e37: x = 16'h3782; 14'h e38: x = 16'h3781; 14'h e39: x = 16'h3780; 14'h e3a: x = 16'h377e; 14'h e3b: x = 16'h377d; 14'h e3c: x = 16'h377c; 14'h e3d: x = 16'h377a; 14'h e3e: x = 16'h3779; 14'h e3f: x = 16'h3778; 14'h e40: x = 16'h3777; 14'h e41: x = 16'h3775; 14'h e42: x = 16'h3774; 14'h e43: x = 16'h3773; 14'h e44: x = 16'h3771; 14'h e45: x = 16'h3770; 14'h e46: x = 16'h376f; 14'h e47: x = 16'h376d; 14'h e48: x = 16'h376c; 14'h e49: x = 16'h376b; 14'h e4a: x = 16'h376a; 14'h e4b: x = 16'h3768; 14'h e4c: x = 16'h3767; 14'h e4d: x = 16'h3766; 14'h e4e: x = 16'h3764; 14'h e4f: x = 16'h3763; 14'h e50: x = 16'h3762; 14'h e51: x = 16'h3761; 14'h e52: x = 16'h375f; 14'h e53: x = 16'h375e; 14'h e54: x = 16'h375d; 14'h e55: x = 16'h375b; 14'h e56: x = 16'h375a; 14'h e57: x = 16'h3759; 14'h e58: x = 16'h3757; 14'h e59: x = 16'h3756; 14'h e5a: x = 16'h3755; 14'h e5b: x = 16'h3754; 14'h e5c: x = 16'h3752; 14'h e5d: x = 16'h3751; 14'h e5e: x = 16'h3750; 14'h e5f: x = 16'h374e; 14'h e60: x = 16'h374d; 14'h e61: x = 16'h374c; 14'h e62: x = 16'h374b; 14'h e63: x = 16'h3749; 14'h e64: x = 16'h3748; 14'h e65: x = 16'h3747; 14'h e66: x = 16'h3745; 14'h e67: x = 16'h3744; 14'h e68: x = 16'h3743; 14'h e69: x = 16'h3742; 14'h e6a: x = 16'h3740; 14'h e6b: x = 16'h373f; 14'h e6c: x = 16'h373e; 14'h e6d: x = 16'h373c; 14'h e6e: x = 16'h373b; 14'h e6f: x = 16'h373a; 14'h e70: x = 16'h3739; 14'h e71: x = 16'h3737; 14'h e72: x = 16'h3736; 14'h e73: x = 16'h3735; 14'h e74: x = 16'h3733; 14'h e75: x = 16'h3732; 14'h e76: x = 16'h3731; 14'h e77: x = 16'h3730; 14'h e78: x = 16'h372e; 14'h e79: x = 16'h372d; 14'h e7a: x = 16'h372c; 14'h e7b: x = 16'h372a; 14'h e7c: x = 16'h3729; 14'h e7d: x = 16'h3728; 14'h e7e: x = 16'h3727; 14'h e7f: x = 16'h3725; 14'h e80: x = 16'h3724; 14'h e81: x = 16'h3723; 14'h e82: x = 16'h3722; 14'h e83: x = 16'h3720; 14'h e84: x = 16'h371f; 14'h e85: x = 16'h371e; 14'h e86: x = 16'h371c; 14'h e87: x = 16'h371b; 14'h e88: x = 16'h371a; 14'h e89: x = 16'h3719; 14'h e8a: x = 16'h3717; 14'h e8b: x = 16'h3716; 14'h e8c: x = 16'h3715; 14'h e8d: x = 16'h3713; 14'h e8e: x = 16'h3712; 14'h e8f: x = 16'h3711; 14'h e90: x = 16'h3710; 14'h e91: x = 16'h370e; 14'h e92: x = 16'h370d; 14'h e93: x = 16'h370c; 14'h e94: x = 16'h370b; 14'h e95: x = 16'h3709; 14'h e96: x = 16'h3708; 14'h e97: x = 16'h3707; 14'h e98: x = 16'h3705; 14'h e99: x = 16'h3704; 14'h e9a: x = 16'h3703; 14'h e9b: x = 16'h3702; 14'h e9c: x = 16'h3700; 14'h e9d: x = 16'h36ff; 14'h e9e: x = 16'h36fe; 14'h e9f: x = 16'h36fc; 14'h ea0: x = 16'h36fb; 14'h ea1: x = 16'h36fa; 14'h ea2: x = 16'h36f9; 14'h ea3: x = 16'h36f7; 14'h ea4: x = 16'h36f6; 14'h ea5: x = 16'h36f5; 14'h ea6: x = 16'h36f4; 14'h ea7: x = 16'h36f2; 14'h ea8: x = 16'h36f1; 14'h ea9: x = 16'h36f0; 14'h eaa: x = 16'h36ee; 14'h eab: x = 16'h36ed; 14'h eac: x = 16'h36ec; 14'h ead: x = 16'h36eb; 14'h eae: x = 16'h36e9; 14'h eaf: x = 16'h36e8; 14'h eb0: x = 16'h36e7; 14'h eb1: x = 16'h36e6; 14'h eb2: x = 16'h36e4; 14'h eb3: x = 16'h36e3; 14'h eb4: x = 16'h36e2; 14'h eb5: x = 16'h36e1; 14'h eb6: x = 16'h36df; 14'h eb7: x = 16'h36de; 14'h eb8: x = 16'h36dd; 14'h eb9: x = 16'h36db; 14'h eba: x = 16'h36da; 14'h ebb: x = 16'h36d9; 14'h ebc: x = 16'h36d8; 14'h ebd: x = 16'h36d6; 14'h ebe: x = 16'h36d5; 14'h ebf: x = 16'h36d4; 14'h ec0: x = 16'h36d3; 14'h ec1: x = 16'h36d1; 14'h ec2: x = 16'h36d0; 14'h ec3: x = 16'h36cf; 14'h ec4: x = 16'h36ce; 14'h ec5: x = 16'h36cc; 14'h ec6: x = 16'h36cb; 14'h ec7: x = 16'h36ca; 14'h ec8: x = 16'h36c8; 14'h ec9: x = 16'h36c7; 14'h eca: x = 16'h36c6; 14'h ecb: x = 16'h36c5; 14'h ecc: x = 16'h36c3; 14'h ecd: x = 16'h36c2; 14'h ece: x = 16'h36c1; 14'h ecf: x = 16'h36c0; 14'h ed0: x = 16'h36be; 14'h ed1: x = 16'h36bd; 14'h ed2: x = 16'h36bc; 14'h ed3: x = 16'h36bb; 14'h ed4: x = 16'h36b9; 14'h ed5: x = 16'h36b8; 14'h ed6: x = 16'h36b7; 14'h ed7: x = 16'h36b6; 14'h ed8: x = 16'h36b4; 14'h ed9: x = 16'h36b3; 14'h eda: x = 16'h36b2; 14'h edb: x = 16'h36b0; 14'h edc: x = 16'h36af; 14'h edd: x = 16'h36ae; 14'h ede: x = 16'h36ad; 14'h edf: x = 16'h36ab; 14'h ee0: x = 16'h36aa; 14'h ee1: x = 16'h36a9; 14'h ee2: x = 16'h36a8; 14'h ee3: x = 16'h36a6; 14'h ee4: x = 16'h36a5; 14'h ee5: x = 16'h36a4; 14'h ee6: x = 16'h36a3; 14'h ee7: x = 16'h36a1; 14'h ee8: x = 16'h36a0; 14'h ee9: x = 16'h369f; 14'h eea: x = 16'h369e; 14'h eeb: x = 16'h369c; 14'h eec: x = 16'h369b; 14'h eed: x = 16'h369a; 14'h eee: x = 16'h3699; 14'h eef: x = 16'h3697; 14'h ef0: x = 16'h3696; 14'h ef1: x = 16'h3695; 14'h ef2: x = 16'h3694; 14'h ef3: x = 16'h3692; 14'h ef4: x = 16'h3691; 14'h ef5: x = 16'h3690; 14'h ef6: x = 16'h368f; 14'h ef7: x = 16'h368d; 14'h ef8: x = 16'h368c; 14'h ef9: x = 16'h368b; 14'h efa: x = 16'h3689; 14'h efb: x = 16'h3688; 14'h efc: x = 16'h3687; 14'h efd: x = 16'h3686; 14'h efe: x = 16'h3684; 14'h eff: x = 16'h3683; 14'h f00: x = 16'h3682; 14'h f01: x = 16'h3681; 14'h f02: x = 16'h367f; 14'h f03: x = 16'h367e; 14'h f04: x = 16'h367d; 14'h f05: x = 16'h367c; 14'h f06: x = 16'h367a; 14'h f07: x = 16'h3679; 14'h f08: x = 16'h3678; 14'h f09: x = 16'h3677; 14'h f0a: x = 16'h3675; 14'h f0b: x = 16'h3674; 14'h f0c: x = 16'h3673; 14'h f0d: x = 16'h3672; 14'h f0e: x = 16'h3670; 14'h f0f: x = 16'h366f; 14'h f10: x = 16'h366e; 14'h f11: x = 16'h366d; 14'h f12: x = 16'h366b; 14'h f13: x = 16'h366a; 14'h f14: x = 16'h3669; 14'h f15: x = 16'h3668; 14'h f16: x = 16'h3666; 14'h f17: x = 16'h3665; 14'h f18: x = 16'h3664; 14'h f19: x = 16'h3663; 14'h f1a: x = 16'h3661; 14'h f1b: x = 16'h3660; 14'h f1c: x = 16'h365f; 14'h f1d: x = 16'h365e; 14'h f1e: x = 16'h365d; 14'h f1f: x = 16'h365b; 14'h f20: x = 16'h365a; 14'h f21: x = 16'h3659; 14'h f22: x = 16'h3658; 14'h f23: x = 16'h3656; 14'h f24: x = 16'h3655; 14'h f25: x = 16'h3654; 14'h f26: x = 16'h3653; 14'h f27: x = 16'h3651; 14'h f28: x = 16'h3650; 14'h f29: x = 16'h364f; 14'h f2a: x = 16'h364e; 14'h f2b: x = 16'h364c; 14'h f2c: x = 16'h364b; 14'h f2d: x = 16'h364a; 14'h f2e: x = 16'h3649; 14'h f2f: x = 16'h3647; 14'h f30: x = 16'h3646; 14'h f31: x = 16'h3645; 14'h f32: x = 16'h3644; 14'h f33: x = 16'h3642; 14'h f34: x = 16'h3641; 14'h f35: x = 16'h3640; 14'h f36: x = 16'h363f; 14'h f37: x = 16'h363d; 14'h f38: x = 16'h363c; 14'h f39: x = 16'h363b; 14'h f3a: x = 16'h363a; 14'h f3b: x = 16'h3638; 14'h f3c: x = 16'h3637; 14'h f3d: x = 16'h3636; 14'h f3e: x = 16'h3635; 14'h f3f: x = 16'h3633; 14'h f40: x = 16'h3632; 14'h f41: x = 16'h3631; 14'h f42: x = 16'h3630; 14'h f43: x = 16'h362f; 14'h f44: x = 16'h362d; 14'h f45: x = 16'h362c; 14'h f46: x = 16'h362b; 14'h f47: x = 16'h362a; 14'h f48: x = 16'h3628; 14'h f49: x = 16'h3627; 14'h f4a: x = 16'h3626; 14'h f4b: x = 16'h3625; 14'h f4c: x = 16'h3623; 14'h f4d: x = 16'h3622; 14'h f4e: x = 16'h3621; 14'h f4f: x = 16'h3620; 14'h f50: x = 16'h361e; 14'h f51: x = 16'h361d; 14'h f52: x = 16'h361c; 14'h f53: x = 16'h361b; 14'h f54: x = 16'h361a; 14'h f55: x = 16'h3618; 14'h f56: x = 16'h3617; 14'h f57: x = 16'h3616; 14'h f58: x = 16'h3615; 14'h f59: x = 16'h3613; 14'h f5a: x = 16'h3612; 14'h f5b: x = 16'h3611; 14'h f5c: x = 16'h3610; 14'h f5d: x = 16'h360e; 14'h f5e: x = 16'h360d; 14'h f5f: x = 16'h360c; 14'h f60: x = 16'h360b; 14'h f61: x = 16'h3609; 14'h f62: x = 16'h3608; 14'h f63: x = 16'h3607; 14'h f64: x = 16'h3606; 14'h f65: x = 16'h3605; 14'h f66: x = 16'h3603; 14'h f67: x = 16'h3602; 14'h f68: x = 16'h3601; 14'h f69: x = 16'h3600; 14'h f6a: x = 16'h35fe; 14'h f6b: x = 16'h35fd; 14'h f6c: x = 16'h35fc; 14'h f6d: x = 16'h35fb; 14'h f6e: x = 16'h35f9; 14'h f6f: x = 16'h35f8; 14'h f70: x = 16'h35f7; 14'h f71: x = 16'h35f6; 14'h f72: x = 16'h35f5; 14'h f73: x = 16'h35f3; 14'h f74: x = 16'h35f2; 14'h f75: x = 16'h35f1; 14'h f76: x = 16'h35f0; 14'h f77: x = 16'h35ee; 14'h f78: x = 16'h35ed; 14'h f79: x = 16'h35ec; 14'h f7a: x = 16'h35eb; 14'h f7b: x = 16'h35ea; 14'h f7c: x = 16'h35e8; 14'h f7d: x = 16'h35e7; 14'h f7e: x = 16'h35e6; 14'h f7f: x = 16'h35e5; 14'h f80: x = 16'h35e3; 14'h f81: x = 16'h35e2; 14'h f82: x = 16'h35e1; 14'h f83: x = 16'h35e0; 14'h f84: x = 16'h35de; 14'h f85: x = 16'h35dd; 14'h f86: x = 16'h35dc; 14'h f87: x = 16'h35db; 14'h f88: x = 16'h35da; 14'h f89: x = 16'h35d8; 14'h f8a: x = 16'h35d7; 14'h f8b: x = 16'h35d6; 14'h f8c: x = 16'h35d5; 14'h f8d: x = 16'h35d3; 14'h f8e: x = 16'h35d2; 14'h f8f: x = 16'h35d1; 14'h f90: x = 16'h35d0; 14'h f91: x = 16'h35cf; 14'h f92: x = 16'h35cd; 14'h f93: x = 16'h35cc; 14'h f94: x = 16'h35cb; 14'h f95: x = 16'h35ca; 14'h f96: x = 16'h35c8; 14'h f97: x = 16'h35c7; 14'h f98: x = 16'h35c6; 14'h f99: x = 16'h35c5; 14'h f9a: x = 16'h35c4; 14'h f9b: x = 16'h35c2; 14'h f9c: x = 16'h35c1; 14'h f9d: x = 16'h35c0; 14'h f9e: x = 16'h35bf; 14'h f9f: x = 16'h35bd; 14'h fa0: x = 16'h35bc; 14'h fa1: x = 16'h35bb; 14'h fa2: x = 16'h35ba; 14'h fa3: x = 16'h35b9; 14'h fa4: x = 16'h35b7; 14'h fa5: x = 16'h35b6; 14'h fa6: x = 16'h35b5; 14'h fa7: x = 16'h35b4; 14'h fa8: x = 16'h35b3; 14'h fa9: x = 16'h35b1; 14'h faa: x = 16'h35b0; 14'h fab: x = 16'h35af; 14'h fac: x = 16'h35ae; 14'h fad: x = 16'h35ac; 14'h fae: x = 16'h35ab; 14'h faf: x = 16'h35aa; 14'h fb0: x = 16'h35a9; 14'h fb1: x = 16'h35a8; 14'h fb2: x = 16'h35a6; 14'h fb3: x = 16'h35a5; 14'h fb4: x = 16'h35a4; 14'h fb5: x = 16'h35a3; 14'h fb6: x = 16'h35a1; 14'h fb7: x = 16'h35a0; 14'h fb8: x = 16'h359f; 14'h fb9: x = 16'h359e; 14'h fba: x = 16'h359d; 14'h fbb: x = 16'h359b; 14'h fbc: x = 16'h359a; 14'h fbd: x = 16'h3599; 14'h fbe: x = 16'h3598; 14'h fbf: x = 16'h3597; 14'h fc0: x = 16'h3595; 14'h fc1: x = 16'h3594; 14'h fc2: x = 16'h3593; 14'h fc3: x = 16'h3592; 14'h fc4: x = 16'h3590; 14'h fc5: x = 16'h358f; 14'h fc6: x = 16'h358e; 14'h fc7: x = 16'h358d; 14'h fc8: x = 16'h358c; 14'h fc9: x = 16'h358a; 14'h fca: x = 16'h3589; 14'h fcb: x = 16'h3588; 14'h fcc: x = 16'h3587; 14'h fcd: x = 16'h3586; 14'h fce: x = 16'h3584; 14'h fcf: x = 16'h3583; 14'h fd0: x = 16'h3582; 14'h fd1: x = 16'h3581; 14'h fd2: x = 16'h3580; 14'h fd3: x = 16'h357e; 14'h fd4: x = 16'h357d; 14'h fd5: x = 16'h357c; 14'h fd6: x = 16'h357b; 14'h fd7: x = 16'h3579; 14'h fd8: x = 16'h3578; 14'h fd9: x = 16'h3577; 14'h fda: x = 16'h3576; 14'h fdb: x = 16'h3575; 14'h fdc: x = 16'h3573; 14'h fdd: x = 16'h3572; 14'h fde: x = 16'h3571; 14'h fdf: x = 16'h3570; 14'h fe0: x = 16'h356f; 14'h fe1: x = 16'h356d; 14'h fe2: x = 16'h356c; 14'h fe3: x = 16'h356b; 14'h fe4: x = 16'h356a; 14'h fe5: x = 16'h3569; 14'h fe6: x = 16'h3567; 14'h fe7: x = 16'h3566; 14'h fe8: x = 16'h3565; 14'h fe9: x = 16'h3564; 14'h fea: x = 16'h3563; 14'h feb: x = 16'h3561; 14'h fec: x = 16'h3560; 14'h fed: x = 16'h355f; 14'h fee: x = 16'h355e; 14'h fef: x = 16'h355d; 14'h ff0: x = 16'h355b; 14'h ff1: x = 16'h355a; 14'h ff2: x = 16'h3559; 14'h ff3: x = 16'h3558; 14'h ff4: x = 16'h3557; 14'h ff5: x = 16'h3555; 14'h ff6: x = 16'h3554; 14'h ff7: x = 16'h3553; 14'h ff8: x = 16'h3552; 14'h ff9: x = 16'h3550; 14'h ffa: x = 16'h354f; 14'h ffb: x = 16'h354e; 14'h ffc: x = 16'h354d; 14'h ffd: x = 16'h354c; 14'h ffe: x = 16'h354a; 14'h fff: x = 16'h3549; 14'h1000: x = 16'h3548; 14'h1001: x = 16'h3547; 14'h1002: x = 16'h3546; 14'h1003: x = 16'h3544; 14'h1004: x = 16'h3543; 14'h1005: x = 16'h3542; 14'h1006: x = 16'h3541; 14'h1007: x = 16'h3540; 14'h1008: x = 16'h353e; 14'h1009: x = 16'h353d; 14'h100a: x = 16'h353c; 14'h100b: x = 16'h353b; 14'h100c: x = 16'h353a; 14'h100d: x = 16'h3538; 14'h100e: x = 16'h3537; 14'h100f: x = 16'h3536; 14'h1010: x = 16'h3535; 14'h1011: x = 16'h3534; 14'h1012: x = 16'h3532; 14'h1013: x = 16'h3531; 14'h1014: x = 16'h3530; 14'h1015: x = 16'h352f; 14'h1016: x = 16'h352e; 14'h1017: x = 16'h352c; 14'h1018: x = 16'h352b; 14'h1019: x = 16'h352a; 14'h101a: x = 16'h3529; 14'h101b: x = 16'h3528; 14'h101c: x = 16'h3527; 14'h101d: x = 16'h3525; 14'h101e: x = 16'h3524; 14'h101f: x = 16'h3523; 14'h1020: x = 16'h3522; 14'h1021: x = 16'h3521; 14'h1022: x = 16'h351f; 14'h1023: x = 16'h351e; 14'h1024: x = 16'h351d; 14'h1025: x = 16'h351c; 14'h1026: x = 16'h351b; 14'h1027: x = 16'h3519; 14'h1028: x = 16'h3518; 14'h1029: x = 16'h3517; 14'h102a: x = 16'h3516; 14'h102b: x = 16'h3515; 14'h102c: x = 16'h3513; 14'h102d: x = 16'h3512; 14'h102e: x = 16'h3511; 14'h102f: x = 16'h3510; 14'h1030: x = 16'h350f; 14'h1031: x = 16'h350d; 14'h1032: x = 16'h350c; 14'h1033: x = 16'h350b; 14'h1034: x = 16'h350a; 14'h1035: x = 16'h3509; 14'h1036: x = 16'h3507; 14'h1037: x = 16'h3506; 14'h1038: x = 16'h3505; 14'h1039: x = 16'h3504; 14'h103a: x = 16'h3503; 14'h103b: x = 16'h3502; 14'h103c: x = 16'h3500; 14'h103d: x = 16'h34ff; 14'h103e: x = 16'h34fe; 14'h103f: x = 16'h34fd; 14'h1040: x = 16'h34fc; 14'h1041: x = 16'h34fa; 14'h1042: x = 16'h34f9; 14'h1043: x = 16'h34f8; 14'h1044: x = 16'h34f7; 14'h1045: x = 16'h34f6; 14'h1046: x = 16'h34f4; 14'h1047: x = 16'h34f3; 14'h1048: x = 16'h34f2; 14'h1049: x = 16'h34f1; 14'h104a: x = 16'h34f0; 14'h104b: x = 16'h34ef; 14'h104c: x = 16'h34ed; 14'h104d: x = 16'h34ec; 14'h104e: x = 16'h34eb; 14'h104f: x = 16'h34ea; 14'h1050: x = 16'h34e9; 14'h1051: x = 16'h34e7; 14'h1052: x = 16'h34e6; 14'h1053: x = 16'h34e5; 14'h1054: x = 16'h34e4; 14'h1055: x = 16'h34e3; 14'h1056: x = 16'h34e1; 14'h1057: x = 16'h34e0; 14'h1058: x = 16'h34df; 14'h1059: x = 16'h34de; 14'h105a: x = 16'h34dd; 14'h105b: x = 16'h34dc; 14'h105c: x = 16'h34da; 14'h105d: x = 16'h34d9; 14'h105e: x = 16'h34d8; 14'h105f: x = 16'h34d7; 14'h1060: x = 16'h34d6; 14'h1061: x = 16'h34d4; 14'h1062: x = 16'h34d3; 14'h1063: x = 16'h34d2; 14'h1064: x = 16'h34d1; 14'h1065: x = 16'h34d0; 14'h1066: x = 16'h34cf; 14'h1067: x = 16'h34cd; 14'h1068: x = 16'h34cc; 14'h1069: x = 16'h34cb; 14'h106a: x = 16'h34ca; 14'h106b: x = 16'h34c9; 14'h106c: x = 16'h34c7; 14'h106d: x = 16'h34c6; 14'h106e: x = 16'h34c5; 14'h106f: x = 16'h34c4; 14'h1070: x = 16'h34c3; 14'h1071: x = 16'h34c2; 14'h1072: x = 16'h34c0; 14'h1073: x = 16'h34bf; 14'h1074: x = 16'h34be; 14'h1075: x = 16'h34bd; 14'h1076: x = 16'h34bc; 14'h1077: x = 16'h34ba; 14'h1078: x = 16'h34b9; 14'h1079: x = 16'h34b8; 14'h107a: x = 16'h34b7; 14'h107b: x = 16'h34b6; 14'h107c: x = 16'h34b5; 14'h107d: x = 16'h34b3; 14'h107e: x = 16'h34b2; 14'h107f: x = 16'h34b1; 14'h1080: x = 16'h34b0; 14'h1081: x = 16'h34af; 14'h1082: x = 16'h34ad; 14'h1083: x = 16'h34ac; 14'h1084: x = 16'h34ab; 14'h1085: x = 16'h34aa; 14'h1086: x = 16'h34a9; 14'h1087: x = 16'h34a8; 14'h1088: x = 16'h34a6; 14'h1089: x = 16'h34a5; 14'h108a: x = 16'h34a4; 14'h108b: x = 16'h34a3; 14'h108c: x = 16'h34a2; 14'h108d: x = 16'h34a1; 14'h108e: x = 16'h349f; 14'h108f: x = 16'h349e; 14'h1090: x = 16'h349d; 14'h1091: x = 16'h349c; 14'h1092: x = 16'h349b; 14'h1093: x = 16'h3499; 14'h1094: x = 16'h3498; 14'h1095: x = 16'h3497; 14'h1096: x = 16'h3496; 14'h1097: x = 16'h3495; 14'h1098: x = 16'h3494; 14'h1099: x = 16'h3492; 14'h109a: x = 16'h3491; 14'h109b: x = 16'h3490; 14'h109c: x = 16'h348f; 14'h109d: x = 16'h348e; 14'h109e: x = 16'h348d; 14'h109f: x = 16'h348b; 14'h10a0: x = 16'h348a; 14'h10a1: x = 16'h3489; 14'h10a2: x = 16'h3488; 14'h10a3: x = 16'h3487; 14'h10a4: x = 16'h3486; 14'h10a5: x = 16'h3484; 14'h10a6: x = 16'h3483; 14'h10a7: x = 16'h3482; 14'h10a8: x = 16'h3481; 14'h10a9: x = 16'h3480; 14'h10aa: x = 16'h347f; 14'h10ab: x = 16'h347d; 14'h10ac: x = 16'h347c; 14'h10ad: x = 16'h347b; 14'h10ae: x = 16'h347a; 14'h10af: x = 16'h3479; 14'h10b0: x = 16'h3477; 14'h10b1: x = 16'h3476; 14'h10b2: x = 16'h3475; 14'h10b3: x = 16'h3474; 14'h10b4: x = 16'h3473; 14'h10b5: x = 16'h3472; 14'h10b6: x = 16'h3470; 14'h10b7: x = 16'h346f; 14'h10b8: x = 16'h346e; 14'h10b9: x = 16'h346d; 14'h10ba: x = 16'h346c; 14'h10bb: x = 16'h346b; 14'h10bc: x = 16'h3469; 14'h10bd: x = 16'h3468; 14'h10be: x = 16'h3467; 14'h10bf: x = 16'h3466; 14'h10c0: x = 16'h3465; 14'h10c1: x = 16'h3464; 14'h10c2: x = 16'h3462; 14'h10c3: x = 16'h3461; 14'h10c4: x = 16'h3460; 14'h10c5: x = 16'h345f; 14'h10c6: x = 16'h345e; 14'h10c7: x = 16'h345d; 14'h10c8: x = 16'h345b; 14'h10c9: x = 16'h345a; 14'h10ca: x = 16'h3459; 14'h10cb: x = 16'h3458; 14'h10cc: x = 16'h3457; 14'h10cd: x = 16'h3456; 14'h10ce: x = 16'h3454; 14'h10cf: x = 16'h3453; 14'h10d0: x = 16'h3452; 14'h10d1: x = 16'h3451; 14'h10d2: x = 16'h3450; 14'h10d3: x = 16'h344f; 14'h10d4: x = 16'h344e; 14'h10d5: x = 16'h344c; 14'h10d6: x = 16'h344b; 14'h10d7: x = 16'h344a; 14'h10d8: x = 16'h3449; 14'h10d9: x = 16'h3448; 14'h10da: x = 16'h3447; 14'h10db: x = 16'h3445; 14'h10dc: x = 16'h3444; 14'h10dd: x = 16'h3443; 14'h10de: x = 16'h3442; 14'h10df: x = 16'h3441; 14'h10e0: x = 16'h3440; 14'h10e1: x = 16'h343e; 14'h10e2: x = 16'h343d; 14'h10e3: x = 16'h343c; 14'h10e4: x = 16'h343b; 14'h10e5: x = 16'h343a; 14'h10e6: x = 16'h3439; 14'h10e7: x = 16'h3437; 14'h10e8: x = 16'h3436; 14'h10e9: x = 16'h3435; 14'h10ea: x = 16'h3434; 14'h10eb: x = 16'h3433; 14'h10ec: x = 16'h3432; 14'h10ed: x = 16'h3430; 14'h10ee: x = 16'h342f; 14'h10ef: x = 16'h342e; 14'h10f0: x = 16'h342d; 14'h10f1: x = 16'h342c; 14'h10f2: x = 16'h342b; 14'h10f3: x = 16'h342a; 14'h10f4: x = 16'h3428; 14'h10f5: x = 16'h3427; 14'h10f6: x = 16'h3426; 14'h10f7: x = 16'h3425; 14'h10f8: x = 16'h3424; 14'h10f9: x = 16'h3423; 14'h10fa: x = 16'h3421; 14'h10fb: x = 16'h3420; 14'h10fc: x = 16'h341f; 14'h10fd: x = 16'h341e; 14'h10fe: x = 16'h341d; 14'h10ff: x = 16'h341c; 14'h1100: x = 16'h341a; 14'h1101: x = 16'h3419; 14'h1102: x = 16'h3418; 14'h1103: x = 16'h3417; 14'h1104: x = 16'h3416; 14'h1105: x = 16'h3415; 14'h1106: x = 16'h3414; 14'h1107: x = 16'h3412; 14'h1108: x = 16'h3411; 14'h1109: x = 16'h3410; 14'h110a: x = 16'h340f; 14'h110b: x = 16'h340e; 14'h110c: x = 16'h340d; 14'h110d: x = 16'h340b; 14'h110e: x = 16'h340a; 14'h110f: x = 16'h3409; 14'h1110: x = 16'h3408; 14'h1111: x = 16'h3407; 14'h1112: x = 16'h3406; 14'h1113: x = 16'h3405; 14'h1114: x = 16'h3403; 14'h1115: x = 16'h3402; 14'h1116: x = 16'h3401; 14'h1117: x = 16'h3400; 14'h1118: x = 16'h33ff; 14'h1119: x = 16'h33fe; 14'h111a: x = 16'h33fc; 14'h111b: x = 16'h33fb; 14'h111c: x = 16'h33fa; 14'h111d: x = 16'h33f9; 14'h111e: x = 16'h33f8; 14'h111f: x = 16'h33f7; 14'h1120: x = 16'h33f6; 14'h1121: x = 16'h33f4; 14'h1122: x = 16'h33f3; 14'h1123: x = 16'h33f2; 14'h1124: x = 16'h33f1; 14'h1125: x = 16'h33f0; 14'h1126: x = 16'h33ef; 14'h1127: x = 16'h33ee; 14'h1128: x = 16'h33ec; 14'h1129: x = 16'h33eb; 14'h112a: x = 16'h33ea; 14'h112b: x = 16'h33e9; 14'h112c: x = 16'h33e8; 14'h112d: x = 16'h33e7; 14'h112e: x = 16'h33e5; 14'h112f: x = 16'h33e4; 14'h1130: x = 16'h33e3; 14'h1131: x = 16'h33e2; 14'h1132: x = 16'h33e1; 14'h1133: x = 16'h33e0; 14'h1134: x = 16'h33df; 14'h1135: x = 16'h33dd; 14'h1136: x = 16'h33dc; 14'h1137: x = 16'h33db; 14'h1138: x = 16'h33da; 14'h1139: x = 16'h33d9; 14'h113a: x = 16'h33d8; 14'h113b: x = 16'h33d7; 14'h113c: x = 16'h33d5; 14'h113d: x = 16'h33d4; 14'h113e: x = 16'h33d3; 14'h113f: x = 16'h33d2; 14'h1140: x = 16'h33d1; 14'h1141: x = 16'h33d0; 14'h1142: x = 16'h33cf; 14'h1143: x = 16'h33cd; 14'h1144: x = 16'h33cc; 14'h1145: x = 16'h33cb; 14'h1146: x = 16'h33ca; 14'h1147: x = 16'h33c9; 14'h1148: x = 16'h33c8; 14'h1149: x = 16'h33c7; 14'h114a: x = 16'h33c5; 14'h114b: x = 16'h33c4; 14'h114c: x = 16'h33c3; 14'h114d: x = 16'h33c2; 14'h114e: x = 16'h33c1; 14'h114f: x = 16'h33c0; 14'h1150: x = 16'h33bf; 14'h1151: x = 16'h33bd; 14'h1152: x = 16'h33bc; 14'h1153: x = 16'h33bb; 14'h1154: x = 16'h33ba; 14'h1155: x = 16'h33b9; 14'h1156: x = 16'h33b8; 14'h1157: x = 16'h33b7; 14'h1158: x = 16'h33b5; 14'h1159: x = 16'h33b4; 14'h115a: x = 16'h33b3; 14'h115b: x = 16'h33b2; 14'h115c: x = 16'h33b1; 14'h115d: x = 16'h33b0; 14'h115e: x = 16'h33af; 14'h115f: x = 16'h33ad; 14'h1160: x = 16'h33ac; 14'h1161: x = 16'h33ab; 14'h1162: x = 16'h33aa; 14'h1163: x = 16'h33a9; 14'h1164: x = 16'h33a8; 14'h1165: x = 16'h33a7; 14'h1166: x = 16'h33a5; 14'h1167: x = 16'h33a4; 14'h1168: x = 16'h33a3; 14'h1169: x = 16'h33a2; 14'h116a: x = 16'h33a1; 14'h116b: x = 16'h33a0; 14'h116c: x = 16'h339f; 14'h116d: x = 16'h339d; 14'h116e: x = 16'h339c; 14'h116f: x = 16'h339b; 14'h1170: x = 16'h339a; 14'h1171: x = 16'h3399; 14'h1172: x = 16'h3398; 14'h1173: x = 16'h3397; 14'h1174: x = 16'h3395; 14'h1175: x = 16'h3394; 14'h1176: x = 16'h3393; 14'h1177: x = 16'h3392; 14'h1178: x = 16'h3391; 14'h1179: x = 16'h3390; 14'h117a: x = 16'h338f; 14'h117b: x = 16'h338e; 14'h117c: x = 16'h338c; 14'h117d: x = 16'h338b; 14'h117e: x = 16'h338a; 14'h117f: x = 16'h3389; 14'h1180: x = 16'h3388; 14'h1181: x = 16'h3387; 14'h1182: x = 16'h3386; 14'h1183: x = 16'h3384; 14'h1184: x = 16'h3383; 14'h1185: x = 16'h3382; 14'h1186: x = 16'h3381; 14'h1187: x = 16'h3380; 14'h1188: x = 16'h337f; 14'h1189: x = 16'h337e; 14'h118a: x = 16'h337c; 14'h118b: x = 16'h337b; 14'h118c: x = 16'h337a; 14'h118d: x = 16'h3379; 14'h118e: x = 16'h3378; 14'h118f: x = 16'h3377; 14'h1190: x = 16'h3376; 14'h1191: x = 16'h3375; 14'h1192: x = 16'h3373; 14'h1193: x = 16'h3372; 14'h1194: x = 16'h3371; 14'h1195: x = 16'h3370; 14'h1196: x = 16'h336f; 14'h1197: x = 16'h336e; 14'h1198: x = 16'h336d; 14'h1199: x = 16'h336b; 14'h119a: x = 16'h336a; 14'h119b: x = 16'h3369; 14'h119c: x = 16'h3368; 14'h119d: x = 16'h3367; 14'h119e: x = 16'h3366; 14'h119f: x = 16'h3365; 14'h11a0: x = 16'h3364; 14'h11a1: x = 16'h3362; 14'h11a2: x = 16'h3361; 14'h11a3: x = 16'h3360; 14'h11a4: x = 16'h335f; 14'h11a5: x = 16'h335e; 14'h11a6: x = 16'h335d; 14'h11a7: x = 16'h335c; 14'h11a8: x = 16'h335b; 14'h11a9: x = 16'h3359; 14'h11aa: x = 16'h3358; 14'h11ab: x = 16'h3357; 14'h11ac: x = 16'h3356; 14'h11ad: x = 16'h3355; 14'h11ae: x = 16'h3354; 14'h11af: x = 16'h3353; 14'h11b0: x = 16'h3352; 14'h11b1: x = 16'h3350; 14'h11b2: x = 16'h334f; 14'h11b3: x = 16'h334e; 14'h11b4: x = 16'h334d; 14'h11b5: x = 16'h334c; 14'h11b6: x = 16'h334b; 14'h11b7: x = 16'h334a; 14'h11b8: x = 16'h3348; 14'h11b9: x = 16'h3347; 14'h11ba: x = 16'h3346; 14'h11bb: x = 16'h3345; 14'h11bc: x = 16'h3344; 14'h11bd: x = 16'h3343; 14'h11be: x = 16'h3342; 14'h11bf: x = 16'h3341; 14'h11c0: x = 16'h333f; 14'h11c1: x = 16'h333e; 14'h11c2: x = 16'h333d; 14'h11c3: x = 16'h333c; 14'h11c4: x = 16'h333b; 14'h11c5: x = 16'h333a; 14'h11c6: x = 16'h3339; 14'h11c7: x = 16'h3338; 14'h11c8: x = 16'h3336; 14'h11c9: x = 16'h3335; 14'h11ca: x = 16'h3334; 14'h11cb: x = 16'h3333; 14'h11cc: x = 16'h3332; 14'h11cd: x = 16'h3331; 14'h11ce: x = 16'h3330; 14'h11cf: x = 16'h332f; 14'h11d0: x = 16'h332d; 14'h11d1: x = 16'h332c; 14'h11d2: x = 16'h332b; 14'h11d3: x = 16'h332a; 14'h11d4: x = 16'h3329; 14'h11d5: x = 16'h3328; 14'h11d6: x = 16'h3327; 14'h11d7: x = 16'h3326; 14'h11d8: x = 16'h3325; 14'h11d9: x = 16'h3323; 14'h11da: x = 16'h3322; 14'h11db: x = 16'h3321; 14'h11dc: x = 16'h3320; 14'h11dd: x = 16'h331f; 14'h11de: x = 16'h331e; 14'h11df: x = 16'h331d; 14'h11e0: x = 16'h331c; 14'h11e1: x = 16'h331a; 14'h11e2: x = 16'h3319; 14'h11e3: x = 16'h3318; 14'h11e4: x = 16'h3317; 14'h11e5: x = 16'h3316; 14'h11e6: x = 16'h3315; 14'h11e7: x = 16'h3314; 14'h11e8: x = 16'h3313; 14'h11e9: x = 16'h3311; 14'h11ea: x = 16'h3310; 14'h11eb: x = 16'h330f; 14'h11ec: x = 16'h330e; 14'h11ed: x = 16'h330d; 14'h11ee: x = 16'h330c; 14'h11ef: x = 16'h330b; 14'h11f0: x = 16'h330a; 14'h11f1: x = 16'h3309; 14'h11f2: x = 16'h3307; 14'h11f3: x = 16'h3306; 14'h11f4: x = 16'h3305; 14'h11f5: x = 16'h3304; 14'h11f6: x = 16'h3303; 14'h11f7: x = 16'h3302; 14'h11f8: x = 16'h3301; 14'h11f9: x = 16'h3300; 14'h11fa: x = 16'h32fe; 14'h11fb: x = 16'h32fd; 14'h11fc: x = 16'h32fc; 14'h11fd: x = 16'h32fb; 14'h11fe: x = 16'h32fa; 14'h11ff: x = 16'h32f9; 14'h1200: x = 16'h32f8; 14'h1201: x = 16'h32f7; 14'h1202: x = 16'h32f6; 14'h1203: x = 16'h32f4; 14'h1204: x = 16'h32f3; 14'h1205: x = 16'h32f2; 14'h1206: x = 16'h32f1; 14'h1207: x = 16'h32f0; 14'h1208: x = 16'h32ef; 14'h1209: x = 16'h32ee; 14'h120a: x = 16'h32ed; 14'h120b: x = 16'h32eb; 14'h120c: x = 16'h32ea; 14'h120d: x = 16'h32e9; 14'h120e: x = 16'h32e8; 14'h120f: x = 16'h32e7; 14'h1210: x = 16'h32e6; 14'h1211: x = 16'h32e5; 14'h1212: x = 16'h32e4; 14'h1213: x = 16'h32e3; 14'h1214: x = 16'h32e1; 14'h1215: x = 16'h32e0; 14'h1216: x = 16'h32df; 14'h1217: x = 16'h32de; 14'h1218: x = 16'h32dd; 14'h1219: x = 16'h32dc; 14'h121a: x = 16'h32db; 14'h121b: x = 16'h32da; 14'h121c: x = 16'h32d9; 14'h121d: x = 16'h32d7; 14'h121e: x = 16'h32d6; 14'h121f: x = 16'h32d5; 14'h1220: x = 16'h32d4; 14'h1221: x = 16'h32d3; 14'h1222: x = 16'h32d2; 14'h1223: x = 16'h32d1; 14'h1224: x = 16'h32d0; 14'h1225: x = 16'h32cf; 14'h1226: x = 16'h32cd; 14'h1227: x = 16'h32cc; 14'h1228: x = 16'h32cb; 14'h1229: x = 16'h32ca; 14'h122a: x = 16'h32c9; 14'h122b: x = 16'h32c8; 14'h122c: x = 16'h32c7; 14'h122d: x = 16'h32c6; 14'h122e: x = 16'h32c5; 14'h122f: x = 16'h32c3; 14'h1230: x = 16'h32c2; 14'h1231: x = 16'h32c1; 14'h1232: x = 16'h32c0; 14'h1233: x = 16'h32bf; 14'h1234: x = 16'h32be; 14'h1235: x = 16'h32bd; 14'h1236: x = 16'h32bc; 14'h1237: x = 16'h32bb; 14'h1238: x = 16'h32b9; 14'h1239: x = 16'h32b8; 14'h123a: x = 16'h32b7; 14'h123b: x = 16'h32b6; 14'h123c: x = 16'h32b5; 14'h123d: x = 16'h32b4; 14'h123e: x = 16'h32b3; 14'h123f: x = 16'h32b2; 14'h1240: x = 16'h32b1; 14'h1241: x = 16'h32b0; 14'h1242: x = 16'h32ae; 14'h1243: x = 16'h32ad; 14'h1244: x = 16'h32ac; 14'h1245: x = 16'h32ab; 14'h1246: x = 16'h32aa; 14'h1247: x = 16'h32a9; 14'h1248: x = 16'h32a8; 14'h1249: x = 16'h32a7; 14'h124a: x = 16'h32a6; 14'h124b: x = 16'h32a4; 14'h124c: x = 16'h32a3; 14'h124d: x = 16'h32a2; 14'h124e: x = 16'h32a1; 14'h124f: x = 16'h32a0; 14'h1250: x = 16'h329f; 14'h1251: x = 16'h329e; 14'h1252: x = 16'h329d; 14'h1253: x = 16'h329c; 14'h1254: x = 16'h329b; 14'h1255: x = 16'h3299; 14'h1256: x = 16'h3298; 14'h1257: x = 16'h3297; 14'h1258: x = 16'h3296; 14'h1259: x = 16'h3295; 14'h125a: x = 16'h3294; 14'h125b: x = 16'h3293; 14'h125c: x = 16'h3292; 14'h125d: x = 16'h3291; 14'h125e: x = 16'h328f; 14'h125f: x = 16'h328e; 14'h1260: x = 16'h328d; 14'h1261: x = 16'h328c; 14'h1262: x = 16'h328b; 14'h1263: x = 16'h328a; 14'h1264: x = 16'h3289; 14'h1265: x = 16'h3288; 14'h1266: x = 16'h3287; 14'h1267: x = 16'h3286; 14'h1268: x = 16'h3284; 14'h1269: x = 16'h3283; 14'h126a: x = 16'h3282; 14'h126b: x = 16'h3281; 14'h126c: x = 16'h3280; 14'h126d: x = 16'h327f; 14'h126e: x = 16'h327e; 14'h126f: x = 16'h327d; 14'h1270: x = 16'h327c; 14'h1271: x = 16'h327b; 14'h1272: x = 16'h3279; 14'h1273: x = 16'h3278; 14'h1274: x = 16'h3277; 14'h1275: x = 16'h3276; 14'h1276: x = 16'h3275; 14'h1277: x = 16'h3274; 14'h1278: x = 16'h3273; 14'h1279: x = 16'h3272; 14'h127a: x = 16'h3271; 14'h127b: x = 16'h3270; 14'h127c: x = 16'h326e; 14'h127d: x = 16'h326d; 14'h127e: x = 16'h326c; 14'h127f: x = 16'h326b; 14'h1280: x = 16'h326a; 14'h1281: x = 16'h3269; 14'h1282: x = 16'h3268; 14'h1283: x = 16'h3267; 14'h1284: x = 16'h3266; 14'h1285: x = 16'h3265; 14'h1286: x = 16'h3263; 14'h1287: x = 16'h3262; 14'h1288: x = 16'h3261; 14'h1289: x = 16'h3260; 14'h128a: x = 16'h325f; 14'h128b: x = 16'h325e; 14'h128c: x = 16'h325d; 14'h128d: x = 16'h325c; 14'h128e: x = 16'h325b; 14'h128f: x = 16'h325a; 14'h1290: x = 16'h3259; 14'h1291: x = 16'h3257; 14'h1292: x = 16'h3256; 14'h1293: x = 16'h3255; 14'h1294: x = 16'h3254; 14'h1295: x = 16'h3253; 14'h1296: x = 16'h3252; 14'h1297: x = 16'h3251; 14'h1298: x = 16'h3250; 14'h1299: x = 16'h324f; 14'h129a: x = 16'h324e; 14'h129b: x = 16'h324c; 14'h129c: x = 16'h324b; 14'h129d: x = 16'h324a; 14'h129e: x = 16'h3249; 14'h129f: x = 16'h3248; 14'h12a0: x = 16'h3247; 14'h12a1: x = 16'h3246; 14'h12a2: x = 16'h3245; 14'h12a3: x = 16'h3244; 14'h12a4: x = 16'h3243; 14'h12a5: x = 16'h3242; 14'h12a6: x = 16'h3240; 14'h12a7: x = 16'h323f; 14'h12a8: x = 16'h323e; 14'h12a9: x = 16'h323d; 14'h12aa: x = 16'h323c; 14'h12ab: x = 16'h323b; 14'h12ac: x = 16'h323a; 14'h12ad: x = 16'h3239; 14'h12ae: x = 16'h3238; 14'h12af: x = 16'h3237; 14'h12b0: x = 16'h3236; 14'h12b1: x = 16'h3234; 14'h12b2: x = 16'h3233; 14'h12b3: x = 16'h3232; 14'h12b4: x = 16'h3231; 14'h12b5: x = 16'h3230; 14'h12b6: x = 16'h322f; 14'h12b7: x = 16'h322e; 14'h12b8: x = 16'h322d; 14'h12b9: x = 16'h322c; 14'h12ba: x = 16'h322b; 14'h12bb: x = 16'h322a; 14'h12bc: x = 16'h3228; 14'h12bd: x = 16'h3227; 14'h12be: x = 16'h3226; 14'h12bf: x = 16'h3225; 14'h12c0: x = 16'h3224; 14'h12c1: x = 16'h3223; 14'h12c2: x = 16'h3222; 14'h12c3: x = 16'h3221; 14'h12c4: x = 16'h3220; 14'h12c5: x = 16'h321f; 14'h12c6: x = 16'h321e; 14'h12c7: x = 16'h321c; 14'h12c8: x = 16'h321b; 14'h12c9: x = 16'h321a; 14'h12ca: x = 16'h3219; 14'h12cb: x = 16'h3218; 14'h12cc: x = 16'h3217; 14'h12cd: x = 16'h3216; 14'h12ce: x = 16'h3215; 14'h12cf: x = 16'h3214; 14'h12d0: x = 16'h3213; 14'h12d1: x = 16'h3212; 14'h12d2: x = 16'h3210; 14'h12d3: x = 16'h320f; 14'h12d4: x = 16'h320e; 14'h12d5: x = 16'h320d; 14'h12d6: x = 16'h320c; 14'h12d7: x = 16'h320b; 14'h12d8: x = 16'h320a; 14'h12d9: x = 16'h3209; 14'h12da: x = 16'h3208; 14'h12db: x = 16'h3207; 14'h12dc: x = 16'h3206; 14'h12dd: x = 16'h3205; 14'h12de: x = 16'h3203; 14'h12df: x = 16'h3202; 14'h12e0: x = 16'h3201; 14'h12e1: x = 16'h3200; 14'h12e2: x = 16'h31ff; 14'h12e3: x = 16'h31fe; 14'h12e4: x = 16'h31fd; 14'h12e5: x = 16'h31fc; 14'h12e6: x = 16'h31fb; 14'h12e7: x = 16'h31fa; 14'h12e8: x = 16'h31f9; 14'h12e9: x = 16'h31f8; 14'h12ea: x = 16'h31f6; 14'h12eb: x = 16'h31f5; 14'h12ec: x = 16'h31f4; 14'h12ed: x = 16'h31f3; 14'h12ee: x = 16'h31f2; 14'h12ef: x = 16'h31f1; 14'h12f0: x = 16'h31f0; 14'h12f1: x = 16'h31ef; 14'h12f2: x = 16'h31ee; 14'h12f3: x = 16'h31ed; 14'h12f4: x = 16'h31ec; 14'h12f5: x = 16'h31eb; 14'h12f6: x = 16'h31e9; 14'h12f7: x = 16'h31e8; 14'h12f8: x = 16'h31e7; 14'h12f9: x = 16'h31e6; 14'h12fa: x = 16'h31e5; 14'h12fb: x = 16'h31e4; 14'h12fc: x = 16'h31e3; 14'h12fd: x = 16'h31e2; 14'h12fe: x = 16'h31e1; 14'h12ff: x = 16'h31e0; 14'h1300: x = 16'h31df; 14'h1301: x = 16'h31de; 14'h1302: x = 16'h31dc; 14'h1303: x = 16'h31db; 14'h1304: x = 16'h31da; 14'h1305: x = 16'h31d9; 14'h1306: x = 16'h31d8; 14'h1307: x = 16'h31d7; 14'h1308: x = 16'h31d6; 14'h1309: x = 16'h31d5; 14'h130a: x = 16'h31d4; 14'h130b: x = 16'h31d3; 14'h130c: x = 16'h31d2; 14'h130d: x = 16'h31d1; 14'h130e: x = 16'h31d0; 14'h130f: x = 16'h31ce; 14'h1310: x = 16'h31cd; 14'h1311: x = 16'h31cc; 14'h1312: x = 16'h31cb; 14'h1313: x = 16'h31ca; 14'h1314: x = 16'h31c9; 14'h1315: x = 16'h31c8; 14'h1316: x = 16'h31c7; 14'h1317: x = 16'h31c6; 14'h1318: x = 16'h31c5; 14'h1319: x = 16'h31c4; 14'h131a: x = 16'h31c3; 14'h131b: x = 16'h31c2; 14'h131c: x = 16'h31c0; 14'h131d: x = 16'h31bf; 14'h131e: x = 16'h31be; 14'h131f: x = 16'h31bd; 14'h1320: x = 16'h31bc; 14'h1321: x = 16'h31bb; 14'h1322: x = 16'h31ba; 14'h1323: x = 16'h31b9; 14'h1324: x = 16'h31b8; 14'h1325: x = 16'h31b7; 14'h1326: x = 16'h31b6; 14'h1327: x = 16'h31b5; 14'h1328: x = 16'h31b4; 14'h1329: x = 16'h31b2; 14'h132a: x = 16'h31b1; 14'h132b: x = 16'h31b0; 14'h132c: x = 16'h31af; 14'h132d: x = 16'h31ae; 14'h132e: x = 16'h31ad; 14'h132f: x = 16'h31ac; 14'h1330: x = 16'h31ab; 14'h1331: x = 16'h31aa; 14'h1332: x = 16'h31a9; 14'h1333: x = 16'h31a8; 14'h1334: x = 16'h31a7; 14'h1335: x = 16'h31a6; 14'h1336: x = 16'h31a4; 14'h1337: x = 16'h31a3; 14'h1338: x = 16'h31a2; 14'h1339: x = 16'h31a1; 14'h133a: x = 16'h31a0; 14'h133b: x = 16'h319f; 14'h133c: x = 16'h319e; 14'h133d: x = 16'h319d; 14'h133e: x = 16'h319c; 14'h133f: x = 16'h319b; 14'h1340: x = 16'h319a; 14'h1341: x = 16'h3199; 14'h1342: x = 16'h3198; 14'h1343: x = 16'h3197; 14'h1344: x = 16'h3195; 14'h1345: x = 16'h3194; 14'h1346: x = 16'h3193; 14'h1347: x = 16'h3192; 14'h1348: x = 16'h3191; 14'h1349: x = 16'h3190; 14'h134a: x = 16'h318f; 14'h134b: x = 16'h318e; 14'h134c: x = 16'h318d; 14'h134d: x = 16'h318c; 14'h134e: x = 16'h318b; 14'h134f: x = 16'h318a; 14'h1350: x = 16'h3189; 14'h1351: x = 16'h3188; 14'h1352: x = 16'h3186; 14'h1353: x = 16'h3185; 14'h1354: x = 16'h3184; 14'h1355: x = 16'h3183; 14'h1356: x = 16'h3182; 14'h1357: x = 16'h3181; 14'h1358: x = 16'h3180; 14'h1359: x = 16'h317f; 14'h135a: x = 16'h317e; 14'h135b: x = 16'h317d; 14'h135c: x = 16'h317c; 14'h135d: x = 16'h317b; 14'h135e: x = 16'h317a; 14'h135f: x = 16'h3179; 14'h1360: x = 16'h3177; 14'h1361: x = 16'h3176; 14'h1362: x = 16'h3175; 14'h1363: x = 16'h3174; 14'h1364: x = 16'h3173; 14'h1365: x = 16'h3172; 14'h1366: x = 16'h3171; 14'h1367: x = 16'h3170; 14'h1368: x = 16'h316f; 14'h1369: x = 16'h316e; 14'h136a: x = 16'h316d; 14'h136b: x = 16'h316c; 14'h136c: x = 16'h316b; 14'h136d: x = 16'h316a; 14'h136e: x = 16'h3169; 14'h136f: x = 16'h3167; 14'h1370: x = 16'h3166; 14'h1371: x = 16'h3165; 14'h1372: x = 16'h3164; 14'h1373: x = 16'h3163; 14'h1374: x = 16'h3162; 14'h1375: x = 16'h3161; 14'h1376: x = 16'h3160; 14'h1377: x = 16'h315f; 14'h1378: x = 16'h315e; 14'h1379: x = 16'h315d; 14'h137a: x = 16'h315c; 14'h137b: x = 16'h315b; 14'h137c: x = 16'h315a; 14'h137d: x = 16'h3159; 14'h137e: x = 16'h3157; 14'h137f: x = 16'h3156; 14'h1380: x = 16'h3155; 14'h1381: x = 16'h3154; 14'h1382: x = 16'h3153; 14'h1383: x = 16'h3152; 14'h1384: x = 16'h3151; 14'h1385: x = 16'h3150; 14'h1386: x = 16'h314f; 14'h1387: x = 16'h314e; 14'h1388: x = 16'h314d; 14'h1389: x = 16'h314c; 14'h138a: x = 16'h314b; 14'h138b: x = 16'h314a; 14'h138c: x = 16'h3149; 14'h138d: x = 16'h3148; 14'h138e: x = 16'h3146; 14'h138f: x = 16'h3145; 14'h1390: x = 16'h3144; 14'h1391: x = 16'h3143; 14'h1392: x = 16'h3142; 14'h1393: x = 16'h3141; 14'h1394: x = 16'h3140; 14'h1395: x = 16'h313f; 14'h1396: x = 16'h313e; 14'h1397: x = 16'h313d; 14'h1398: x = 16'h313c; 14'h1399: x = 16'h313b; 14'h139a: x = 16'h313a; 14'h139b: x = 16'h3139; 14'h139c: x = 16'h3138; 14'h139d: x = 16'h3137; 14'h139e: x = 16'h3135; 14'h139f: x = 16'h3134; 14'h13a0: x = 16'h3133; 14'h13a1: x = 16'h3132; 14'h13a2: x = 16'h3131; 14'h13a3: x = 16'h3130; 14'h13a4: x = 16'h312f; 14'h13a5: x = 16'h312e; 14'h13a6: x = 16'h312d; 14'h13a7: x = 16'h312c; 14'h13a8: x = 16'h312b; 14'h13a9: x = 16'h312a; 14'h13aa: x = 16'h3129; 14'h13ab: x = 16'h3128; 14'h13ac: x = 16'h3127; 14'h13ad: x = 16'h3126; 14'h13ae: x = 16'h3125; 14'h13af: x = 16'h3123; 14'h13b0: x = 16'h3122; 14'h13b1: x = 16'h3121; 14'h13b2: x = 16'h3120; 14'h13b3: x = 16'h311f; 14'h13b4: x = 16'h311e; 14'h13b5: x = 16'h311d; 14'h13b6: x = 16'h311c; 14'h13b7: x = 16'h311b; 14'h13b8: x = 16'h311a; 14'h13b9: x = 16'h3119; 14'h13ba: x = 16'h3118; 14'h13bb: x = 16'h3117; 14'h13bc: x = 16'h3116; 14'h13bd: x = 16'h3115; 14'h13be: x = 16'h3114; 14'h13bf: x = 16'h3113; 14'h13c0: x = 16'h3111; 14'h13c1: x = 16'h3110; 14'h13c2: x = 16'h310f; 14'h13c3: x = 16'h310e; 14'h13c4: x = 16'h310d; 14'h13c5: x = 16'h310c; 14'h13c6: x = 16'h310b; 14'h13c7: x = 16'h310a; 14'h13c8: x = 16'h3109; 14'h13c9: x = 16'h3108; 14'h13ca: x = 16'h3107; 14'h13cb: x = 16'h3106; 14'h13cc: x = 16'h3105; 14'h13cd: x = 16'h3104; 14'h13ce: x = 16'h3103; 14'h13cf: x = 16'h3102; 14'h13d0: x = 16'h3101; 14'h13d1: x = 16'h3100; 14'h13d2: x = 16'h30fe; 14'h13d3: x = 16'h30fd; 14'h13d4: x = 16'h30fc; 14'h13d5: x = 16'h30fb; 14'h13d6: x = 16'h30fa; 14'h13d7: x = 16'h30f9; 14'h13d8: x = 16'h30f8; 14'h13d9: x = 16'h30f7; 14'h13da: x = 16'h30f6; 14'h13db: x = 16'h30f5; 14'h13dc: x = 16'h30f4; 14'h13dd: x = 16'h30f3; 14'h13de: x = 16'h30f2; 14'h13df: x = 16'h30f1; 14'h13e0: x = 16'h30f0; 14'h13e1: x = 16'h30ef; 14'h13e2: x = 16'h30ee; 14'h13e3: x = 16'h30ed; 14'h13e4: x = 16'h30ec; 14'h13e5: x = 16'h30ea; 14'h13e6: x = 16'h30e9; 14'h13e7: x = 16'h30e8; 14'h13e8: x = 16'h30e7; 14'h13e9: x = 16'h30e6; 14'h13ea: x = 16'h30e5; 14'h13eb: x = 16'h30e4; 14'h13ec: x = 16'h30e3; 14'h13ed: x = 16'h30e2; 14'h13ee: x = 16'h30e1; 14'h13ef: x = 16'h30e0; 14'h13f0: x = 16'h30df; 14'h13f1: x = 16'h30de; 14'h13f2: x = 16'h30dd; 14'h13f3: x = 16'h30dc; 14'h13f4: x = 16'h30db; 14'h13f5: x = 16'h30da; 14'h13f6: x = 16'h30d9; 14'h13f7: x = 16'h30d8; 14'h13f8: x = 16'h30d7; 14'h13f9: x = 16'h30d5; 14'h13fa: x = 16'h30d4; 14'h13fb: x = 16'h30d3; 14'h13fc: x = 16'h30d2; 14'h13fd: x = 16'h30d1; 14'h13fe: x = 16'h30d0; 14'h13ff: x = 16'h30cf; 14'h1400: x = 16'h30ce; 14'h1401: x = 16'h30cd; 14'h1402: x = 16'h30cc; 14'h1403: x = 16'h30cb; 14'h1404: x = 16'h30ca; 14'h1405: x = 16'h30c9; 14'h1406: x = 16'h30c8; 14'h1407: x = 16'h30c7; 14'h1408: x = 16'h30c6; 14'h1409: x = 16'h30c5; 14'h140a: x = 16'h30c4; 14'h140b: x = 16'h30c3; 14'h140c: x = 16'h30c2; 14'h140d: x = 16'h30c0; 14'h140e: x = 16'h30bf; 14'h140f: x = 16'h30be; 14'h1410: x = 16'h30bd; 14'h1411: x = 16'h30bc; 14'h1412: x = 16'h30bb; 14'h1413: x = 16'h30ba; 14'h1414: x = 16'h30b9; 14'h1415: x = 16'h30b8; 14'h1416: x = 16'h30b7; 14'h1417: x = 16'h30b6; 14'h1418: x = 16'h30b5; 14'h1419: x = 16'h30b4; 14'h141a: x = 16'h30b3; 14'h141b: x = 16'h30b2; 14'h141c: x = 16'h30b1; 14'h141d: x = 16'h30b0; 14'h141e: x = 16'h30af; 14'h141f: x = 16'h30ae; 14'h1420: x = 16'h30ad; 14'h1421: x = 16'h30ac; 14'h1422: x = 16'h30ab; 14'h1423: x = 16'h30a9; 14'h1424: x = 16'h30a8; 14'h1425: x = 16'h30a7; 14'h1426: x = 16'h30a6; 14'h1427: x = 16'h30a5; 14'h1428: x = 16'h30a4; 14'h1429: x = 16'h30a3; 14'h142a: x = 16'h30a2; 14'h142b: x = 16'h30a1; 14'h142c: x = 16'h30a0; 14'h142d: x = 16'h309f; 14'h142e: x = 16'h309e; 14'h142f: x = 16'h309d; 14'h1430: x = 16'h309c; 14'h1431: x = 16'h309b; 14'h1432: x = 16'h309a; 14'h1433: x = 16'h3099; 14'h1434: x = 16'h3098; 14'h1435: x = 16'h3097; 14'h1436: x = 16'h3096; 14'h1437: x = 16'h3095; 14'h1438: x = 16'h3094; 14'h1439: x = 16'h3093; 14'h143a: x = 16'h3091; 14'h143b: x = 16'h3090; 14'h143c: x = 16'h308f; 14'h143d: x = 16'h308e; 14'h143e: x = 16'h308d; 14'h143f: x = 16'h308c; 14'h1440: x = 16'h308b; 14'h1441: x = 16'h308a; 14'h1442: x = 16'h3089; 14'h1443: x = 16'h3088; 14'h1444: x = 16'h3087; 14'h1445: x = 16'h3086; 14'h1446: x = 16'h3085; 14'h1447: x = 16'h3084; 14'h1448: x = 16'h3083; 14'h1449: x = 16'h3082; 14'h144a: x = 16'h3081; 14'h144b: x = 16'h3080; 14'h144c: x = 16'h307f; 14'h144d: x = 16'h307e; 14'h144e: x = 16'h307d; 14'h144f: x = 16'h307c; 14'h1450: x = 16'h307b; 14'h1451: x = 16'h307a; 14'h1452: x = 16'h3078; 14'h1453: x = 16'h3077; 14'h1454: x = 16'h3076; 14'h1455: x = 16'h3075; 14'h1456: x = 16'h3074; 14'h1457: x = 16'h3073; 14'h1458: x = 16'h3072; 14'h1459: x = 16'h3071; 14'h145a: x = 16'h3070; 14'h145b: x = 16'h306f; 14'h145c: x = 16'h306e; 14'h145d: x = 16'h306d; 14'h145e: x = 16'h306c; 14'h145f: x = 16'h306b; 14'h1460: x = 16'h306a; 14'h1461: x = 16'h3069; 14'h1462: x = 16'h3068; 14'h1463: x = 16'h3067; 14'h1464: x = 16'h3066; 14'h1465: x = 16'h3065; 14'h1466: x = 16'h3064; 14'h1467: x = 16'h3063; 14'h1468: x = 16'h3062; 14'h1469: x = 16'h3061; 14'h146a: x = 16'h3060; 14'h146b: x = 16'h305f; 14'h146c: x = 16'h305d; 14'h146d: x = 16'h305c; 14'h146e: x = 16'h305b; 14'h146f: x = 16'h305a; 14'h1470: x = 16'h3059; 14'h1471: x = 16'h3058; 14'h1472: x = 16'h3057; 14'h1473: x = 16'h3056; 14'h1474: x = 16'h3055; 14'h1475: x = 16'h3054; 14'h1476: x = 16'h3053; 14'h1477: x = 16'h3052; 14'h1478: x = 16'h3051; 14'h1479: x = 16'h3050; 14'h147a: x = 16'h304f; 14'h147b: x = 16'h304e; 14'h147c: x = 16'h304d; 14'h147d: x = 16'h304c; 14'h147e: x = 16'h304b; 14'h147f: x = 16'h304a; 14'h1480: x = 16'h3049; 14'h1481: x = 16'h3048; 14'h1482: x = 16'h3047; 14'h1483: x = 16'h3046; 14'h1484: x = 16'h3045; 14'h1485: x = 16'h3044; 14'h1486: x = 16'h3043; 14'h1487: x = 16'h3042; 14'h1488: x = 16'h3041; 14'h1489: x = 16'h303f; 14'h148a: x = 16'h303e; 14'h148b: x = 16'h303d; 14'h148c: x = 16'h303c; 14'h148d: x = 16'h303b; 14'h148e: x = 16'h303a; 14'h148f: x = 16'h3039; 14'h1490: x = 16'h3038; 14'h1491: x = 16'h3037; 14'h1492: x = 16'h3036; 14'h1493: x = 16'h3035; 14'h1494: x = 16'h3034; 14'h1495: x = 16'h3033; 14'h1496: x = 16'h3032; 14'h1497: x = 16'h3031; 14'h1498: x = 16'h3030; 14'h1499: x = 16'h302f; 14'h149a: x = 16'h302e; 14'h149b: x = 16'h302d; 14'h149c: x = 16'h302c; 14'h149d: x = 16'h302b; 14'h149e: x = 16'h302a; 14'h149f: x = 16'h3029; 14'h14a0: x = 16'h3028; 14'h14a1: x = 16'h3027; 14'h14a2: x = 16'h3026; 14'h14a3: x = 16'h3025; 14'h14a4: x = 16'h3024; 14'h14a5: x = 16'h3023; 14'h14a6: x = 16'h3022; 14'h14a7: x = 16'h3021; 14'h14a8: x = 16'h301f; 14'h14a9: x = 16'h301e; 14'h14aa: x = 16'h301d; 14'h14ab: x = 16'h301c; 14'h14ac: x = 16'h301b; 14'h14ad: x = 16'h301a; 14'h14ae: x = 16'h3019; 14'h14af: x = 16'h3018; 14'h14b0: x = 16'h3017; 14'h14b1: x = 16'h3016; 14'h14b2: x = 16'h3015; 14'h14b3: x = 16'h3014; 14'h14b4: x = 16'h3013; 14'h14b5: x = 16'h3012; 14'h14b6: x = 16'h3011; 14'h14b7: x = 16'h3010; 14'h14b8: x = 16'h300f; 14'h14b9: x = 16'h300e; 14'h14ba: x = 16'h300d; 14'h14bb: x = 16'h300c; 14'h14bc: x = 16'h300b; 14'h14bd: x = 16'h300a; 14'h14be: x = 16'h3009; 14'h14bf: x = 16'h3008; 14'h14c0: x = 16'h3007; 14'h14c1: x = 16'h3006; 14'h14c2: x = 16'h3005; 14'h14c3: x = 16'h3004; 14'h14c4: x = 16'h3003; 14'h14c5: x = 16'h3002; 14'h14c6: x = 16'h3001; 14'h14c7: x = 16'h3000; 14'h14c8: x = 16'h2fff; 14'h14c9: x = 16'h2ffe; 14'h14ca: x = 16'h2ffd; 14'h14cb: x = 16'h2ffc; 14'h14cc: x = 16'h2ffa; 14'h14cd: x = 16'h2ff9; 14'h14ce: x = 16'h2ff8; 14'h14cf: x = 16'h2ff7; 14'h14d0: x = 16'h2ff6; 14'h14d1: x = 16'h2ff5; 14'h14d2: x = 16'h2ff4; 14'h14d3: x = 16'h2ff3; 14'h14d4: x = 16'h2ff2; 14'h14d5: x = 16'h2ff1; 14'h14d6: x = 16'h2ff0; 14'h14d7: x = 16'h2fef; 14'h14d8: x = 16'h2fee; 14'h14d9: x = 16'h2fed; 14'h14da: x = 16'h2fec; 14'h14db: x = 16'h2feb; 14'h14dc: x = 16'h2fea; 14'h14dd: x = 16'h2fe9; 14'h14de: x = 16'h2fe8; 14'h14df: x = 16'h2fe7; 14'h14e0: x = 16'h2fe6; 14'h14e1: x = 16'h2fe5; 14'h14e2: x = 16'h2fe4; 14'h14e3: x = 16'h2fe3; 14'h14e4: x = 16'h2fe2; 14'h14e5: x = 16'h2fe1; 14'h14e6: x = 16'h2fe0; 14'h14e7: x = 16'h2fdf; 14'h14e8: x = 16'h2fde; 14'h14e9: x = 16'h2fdd; 14'h14ea: x = 16'h2fdc; 14'h14eb: x = 16'h2fdb; 14'h14ec: x = 16'h2fda; 14'h14ed: x = 16'h2fd9; 14'h14ee: x = 16'h2fd8; 14'h14ef: x = 16'h2fd7; 14'h14f0: x = 16'h2fd6; 14'h14f1: x = 16'h2fd5; 14'h14f2: x = 16'h2fd4; 14'h14f3: x = 16'h2fd3; 14'h14f4: x = 16'h2fd2; 14'h14f5: x = 16'h2fd0; 14'h14f6: x = 16'h2fcf; 14'h14f7: x = 16'h2fce; 14'h14f8: x = 16'h2fcd; 14'h14f9: x = 16'h2fcc; 14'h14fa: x = 16'h2fcb; 14'h14fb: x = 16'h2fca; 14'h14fc: x = 16'h2fc9; 14'h14fd: x = 16'h2fc8; 14'h14fe: x = 16'h2fc7; 14'h14ff: x = 16'h2fc6; 14'h1500: x = 16'h2fc5; 14'h1501: x = 16'h2fc4; 14'h1502: x = 16'h2fc3; 14'h1503: x = 16'h2fc2; 14'h1504: x = 16'h2fc1; 14'h1505: x = 16'h2fc0; 14'h1506: x = 16'h2fbf; 14'h1507: x = 16'h2fbe; 14'h1508: x = 16'h2fbd; 14'h1509: x = 16'h2fbc; 14'h150a: x = 16'h2fbb; 14'h150b: x = 16'h2fba; 14'h150c: x = 16'h2fb9; 14'h150d: x = 16'h2fb8; 14'h150e: x = 16'h2fb7; 14'h150f: x = 16'h2fb6; 14'h1510: x = 16'h2fb5; 14'h1511: x = 16'h2fb4; 14'h1512: x = 16'h2fb3; 14'h1513: x = 16'h2fb2; 14'h1514: x = 16'h2fb1; 14'h1515: x = 16'h2fb0; 14'h1516: x = 16'h2faf; 14'h1517: x = 16'h2fae; 14'h1518: x = 16'h2fad; 14'h1519: x = 16'h2fac; 14'h151a: x = 16'h2fab; 14'h151b: x = 16'h2faa; 14'h151c: x = 16'h2fa9; 14'h151d: x = 16'h2fa8; 14'h151e: x = 16'h2fa7; 14'h151f: x = 16'h2fa6; 14'h1520: x = 16'h2fa5; 14'h1521: x = 16'h2fa4; 14'h1522: x = 16'h2fa3; 14'h1523: x = 16'h2fa2; 14'h1524: x = 16'h2fa1; 14'h1525: x = 16'h2fa0; 14'h1526: x = 16'h2f9f; 14'h1527: x = 16'h2f9e; 14'h1528: x = 16'h2f9d; 14'h1529: x = 16'h2f9b; 14'h152a: x = 16'h2f9a; 14'h152b: x = 16'h2f99; 14'h152c: x = 16'h2f98; 14'h152d: x = 16'h2f97; 14'h152e: x = 16'h2f96; 14'h152f: x = 16'h2f95; 14'h1530: x = 16'h2f94; 14'h1531: x = 16'h2f93; 14'h1532: x = 16'h2f92; 14'h1533: x = 16'h2f91; 14'h1534: x = 16'h2f90; 14'h1535: x = 16'h2f8f; 14'h1536: x = 16'h2f8e; 14'h1537: x = 16'h2f8d; 14'h1538: x = 16'h2f8c; 14'h1539: x = 16'h2f8b; 14'h153a: x = 16'h2f8a; 14'h153b: x = 16'h2f89; 14'h153c: x = 16'h2f88; 14'h153d: x = 16'h2f87; 14'h153e: x = 16'h2f86; 14'h153f: x = 16'h2f85; 14'h1540: x = 16'h2f84; 14'h1541: x = 16'h2f83; 14'h1542: x = 16'h2f82; 14'h1543: x = 16'h2f81; 14'h1544: x = 16'h2f80; 14'h1545: x = 16'h2f7f; 14'h1546: x = 16'h2f7e; 14'h1547: x = 16'h2f7d; 14'h1548: x = 16'h2f7c; 14'h1549: x = 16'h2f7b; 14'h154a: x = 16'h2f7a; 14'h154b: x = 16'h2f79; 14'h154c: x = 16'h2f78; 14'h154d: x = 16'h2f77; 14'h154e: x = 16'h2f76; 14'h154f: x = 16'h2f75; 14'h1550: x = 16'h2f74; 14'h1551: x = 16'h2f73; 14'h1552: x = 16'h2f72; 14'h1553: x = 16'h2f71; 14'h1554: x = 16'h2f70; 14'h1555: x = 16'h2f6f; 14'h1556: x = 16'h2f6e; 14'h1557: x = 16'h2f6d; 14'h1558: x = 16'h2f6c; 14'h1559: x = 16'h2f6b; 14'h155a: x = 16'h2f6a; 14'h155b: x = 16'h2f69; 14'h155c: x = 16'h2f68; 14'h155d: x = 16'h2f67; 14'h155e: x = 16'h2f66; 14'h155f: x = 16'h2f65; 14'h1560: x = 16'h2f64; 14'h1561: x = 16'h2f63; 14'h1562: x = 16'h2f62; 14'h1563: x = 16'h2f61; 14'h1564: x = 16'h2f60; 14'h1565: x = 16'h2f5f; 14'h1566: x = 16'h2f5e; 14'h1567: x = 16'h2f5d; 14'h1568: x = 16'h2f5c; 14'h1569: x = 16'h2f5b; 14'h156a: x = 16'h2f5a; 14'h156b: x = 16'h2f59; 14'h156c: x = 16'h2f58; 14'h156d: x = 16'h2f57; 14'h156e: x = 16'h2f56; 14'h156f: x = 16'h2f55; 14'h1570: x = 16'h2f54; 14'h1571: x = 16'h2f53; 14'h1572: x = 16'h2f52; 14'h1573: x = 16'h2f51; 14'h1574: x = 16'h2f50; 14'h1575: x = 16'h2f4f; 14'h1576: x = 16'h2f4e; 14'h1577: x = 16'h2f4d; 14'h1578: x = 16'h2f4c; 14'h1579: x = 16'h2f4b; 14'h157a: x = 16'h2f49; 14'h157b: x = 16'h2f48; 14'h157c: x = 16'h2f47; 14'h157d: x = 16'h2f46; 14'h157e: x = 16'h2f45; 14'h157f: x = 16'h2f44; 14'h1580: x = 16'h2f43; 14'h1581: x = 16'h2f42; 14'h1582: x = 16'h2f41; 14'h1583: x = 16'h2f40; 14'h1584: x = 16'h2f3f; 14'h1585: x = 16'h2f3e; 14'h1586: x = 16'h2f3d; 14'h1587: x = 16'h2f3c; 14'h1588: x = 16'h2f3b; 14'h1589: x = 16'h2f3a; 14'h158a: x = 16'h2f39; 14'h158b: x = 16'h2f38; 14'h158c: x = 16'h2f37; 14'h158d: x = 16'h2f36; 14'h158e: x = 16'h2f35; 14'h158f: x = 16'h2f34; 14'h1590: x = 16'h2f33; 14'h1591: x = 16'h2f32; 14'h1592: x = 16'h2f31; 14'h1593: x = 16'h2f30; 14'h1594: x = 16'h2f2f; 14'h1595: x = 16'h2f2e; 14'h1596: x = 16'h2f2d; 14'h1597: x = 16'h2f2c; 14'h1598: x = 16'h2f2b; 14'h1599: x = 16'h2f2a; 14'h159a: x = 16'h2f29; 14'h159b: x = 16'h2f28; 14'h159c: x = 16'h2f27; 14'h159d: x = 16'h2f26; 14'h159e: x = 16'h2f25; 14'h159f: x = 16'h2f24; 14'h15a0: x = 16'h2f23; 14'h15a1: x = 16'h2f22; 14'h15a2: x = 16'h2f21; 14'h15a3: x = 16'h2f20; 14'h15a4: x = 16'h2f1f; 14'h15a5: x = 16'h2f1e; 14'h15a6: x = 16'h2f1d; 14'h15a7: x = 16'h2f1c; 14'h15a8: x = 16'h2f1b; 14'h15a9: x = 16'h2f1a; 14'h15aa: x = 16'h2f19; 14'h15ab: x = 16'h2f18; 14'h15ac: x = 16'h2f17; 14'h15ad: x = 16'h2f16; 14'h15ae: x = 16'h2f15; 14'h15af: x = 16'h2f14; 14'h15b0: x = 16'h2f13; 14'h15b1: x = 16'h2f12; 14'h15b2: x = 16'h2f11; 14'h15b3: x = 16'h2f10; 14'h15b4: x = 16'h2f0f; 14'h15b5: x = 16'h2f0e; 14'h15b6: x = 16'h2f0d; 14'h15b7: x = 16'h2f0c; 14'h15b8: x = 16'h2f0b; 14'h15b9: x = 16'h2f0a; 14'h15ba: x = 16'h2f09; 14'h15bb: x = 16'h2f08; 14'h15bc: x = 16'h2f07; 14'h15bd: x = 16'h2f06; 14'h15be: x = 16'h2f05; 14'h15bf: x = 16'h2f04; 14'h15c0: x = 16'h2f03; 14'h15c1: x = 16'h2f02; 14'h15c2: x = 16'h2f01; 14'h15c3: x = 16'h2f00; 14'h15c4: x = 16'h2eff; 14'h15c5: x = 16'h2efe; 14'h15c6: x = 16'h2efd; 14'h15c7: x = 16'h2efc; 14'h15c8: x = 16'h2efb; 14'h15c9: x = 16'h2efa; 14'h15ca: x = 16'h2ef9; 14'h15cb: x = 16'h2ef8; 14'h15cc: x = 16'h2ef7; 14'h15cd: x = 16'h2ef6; 14'h15ce: x = 16'h2ef5; 14'h15cf: x = 16'h2ef4; 14'h15d0: x = 16'h2ef3; 14'h15d1: x = 16'h2ef2; 14'h15d2: x = 16'h2ef1; 14'h15d3: x = 16'h2ef0; 14'h15d4: x = 16'h2eef; 14'h15d5: x = 16'h2eee; 14'h15d6: x = 16'h2eed; 14'h15d7: x = 16'h2eec; 14'h15d8: x = 16'h2eeb; 14'h15d9: x = 16'h2eea; 14'h15da: x = 16'h2ee9; 14'h15db: x = 16'h2ee8; 14'h15dc: x = 16'h2ee7; 14'h15dd: x = 16'h2ee6; 14'h15de: x = 16'h2ee5; 14'h15df: x = 16'h2ee4; 14'h15e0: x = 16'h2ee3; 14'h15e1: x = 16'h2ee2; 14'h15e2: x = 16'h2ee1; 14'h15e3: x = 16'h2ee0; 14'h15e4: x = 16'h2edf; 14'h15e5: x = 16'h2ede; 14'h15e6: x = 16'h2edd; 14'h15e7: x = 16'h2edc; 14'h15e8: x = 16'h2edb; 14'h15e9: x = 16'h2eda; 14'h15ea: x = 16'h2ed9; 14'h15eb: x = 16'h2ed8; 14'h15ec: x = 16'h2ed7; 14'h15ed: x = 16'h2ed6; 14'h15ee: x = 16'h2ed5; 14'h15ef: x = 16'h2ed4; 14'h15f0: x = 16'h2ed3; 14'h15f1: x = 16'h2ed2; 14'h15f2: x = 16'h2ed1; 14'h15f3: x = 16'h2ed0; 14'h15f4: x = 16'h2ecf; 14'h15f5: x = 16'h2ece; 14'h15f6: x = 16'h2ecd; 14'h15f7: x = 16'h2ecc; 14'h15f8: x = 16'h2ecb; 14'h15f9: x = 16'h2eca; 14'h15fa: x = 16'h2ec9; 14'h15fb: x = 16'h2ec8; 14'h15fc: x = 16'h2ec7; 14'h15fd: x = 16'h2ec6; 14'h15fe: x = 16'h2ec5; 14'h15ff: x = 16'h2ec4; 14'h1600: x = 16'h2ec3; 14'h1601: x = 16'h2ec2; 14'h1602: x = 16'h2ec1; 14'h1603: x = 16'h2ec0; 14'h1604: x = 16'h2ebf; 14'h1605: x = 16'h2ebe; 14'h1606: x = 16'h2ebd; 14'h1607: x = 16'h2ebc; 14'h1608: x = 16'h2ebb; 14'h1609: x = 16'h2eba; 14'h160a: x = 16'h2eb9; 14'h160b: x = 16'h2eb8; 14'h160c: x = 16'h2eb7; 14'h160d: x = 16'h2eb6; 14'h160e: x = 16'h2eb5; 14'h160f: x = 16'h2eb4; 14'h1610: x = 16'h2eb3; 14'h1611: x = 16'h2eb2; 14'h1612: x = 16'h2eb1; 14'h1613: x = 16'h2eb0; 14'h1614: x = 16'h2eaf; 14'h1615: x = 16'h2eae; 14'h1616: x = 16'h2ead; 14'h1617: x = 16'h2eac; 14'h1618: x = 16'h2eab; 14'h1619: x = 16'h2eaa; 14'h161a: x = 16'h2ea9; 14'h161b: x = 16'h2ea8; 14'h161c: x = 16'h2ea7; 14'h161d: x = 16'h2ea6; 14'h161e: x = 16'h2ea5; 14'h161f: x = 16'h2ea4; 14'h1620: x = 16'h2ea3; 14'h1621: x = 16'h2ea2; 14'h1622: x = 16'h2ea1; 14'h1623: x = 16'h2ea0; 14'h1624: x = 16'h2e9f; 14'h1625: x = 16'h2e9f; 14'h1626: x = 16'h2e9e; 14'h1627: x = 16'h2e9d; 14'h1628: x = 16'h2e9c; 14'h1629: x = 16'h2e9b; 14'h162a: x = 16'h2e9a; 14'h162b: x = 16'h2e99; 14'h162c: x = 16'h2e98; 14'h162d: x = 16'h2e97; 14'h162e: x = 16'h2e96; 14'h162f: x = 16'h2e95; 14'h1630: x = 16'h2e94; 14'h1631: x = 16'h2e93; 14'h1632: x = 16'h2e92; 14'h1633: x = 16'h2e91; 14'h1634: x = 16'h2e90; 14'h1635: x = 16'h2e8f; 14'h1636: x = 16'h2e8e; 14'h1637: x = 16'h2e8d; 14'h1638: x = 16'h2e8c; 14'h1639: x = 16'h2e8b; 14'h163a: x = 16'h2e8a; 14'h163b: x = 16'h2e89; 14'h163c: x = 16'h2e88; 14'h163d: x = 16'h2e87; 14'h163e: x = 16'h2e86; 14'h163f: x = 16'h2e85; 14'h1640: x = 16'h2e84; 14'h1641: x = 16'h2e83; 14'h1642: x = 16'h2e82; 14'h1643: x = 16'h2e81; 14'h1644: x = 16'h2e80; 14'h1645: x = 16'h2e7f; 14'h1646: x = 16'h2e7e; 14'h1647: x = 16'h2e7d; 14'h1648: x = 16'h2e7c; 14'h1649: x = 16'h2e7b; 14'h164a: x = 16'h2e7a; 14'h164b: x = 16'h2e79; 14'h164c: x = 16'h2e78; 14'h164d: x = 16'h2e77; 14'h164e: x = 16'h2e76; 14'h164f: x = 16'h2e75; 14'h1650: x = 16'h2e74; 14'h1651: x = 16'h2e73; 14'h1652: x = 16'h2e72; 14'h1653: x = 16'h2e71; 14'h1654: x = 16'h2e70; 14'h1655: x = 16'h2e6f; 14'h1656: x = 16'h2e6e; 14'h1657: x = 16'h2e6d; 14'h1658: x = 16'h2e6c; 14'h1659: x = 16'h2e6b; 14'h165a: x = 16'h2e6a; 14'h165b: x = 16'h2e69; 14'h165c: x = 16'h2e68; 14'h165d: x = 16'h2e67; 14'h165e: x = 16'h2e66; 14'h165f: x = 16'h2e65; 14'h1660: x = 16'h2e64; 14'h1661: x = 16'h2e63; 14'h1662: x = 16'h2e62; 14'h1663: x = 16'h2e61; 14'h1664: x = 16'h2e60; 14'h1665: x = 16'h2e5f; 14'h1666: x = 16'h2e5e; 14'h1667: x = 16'h2e5d; 14'h1668: x = 16'h2e5c; 14'h1669: x = 16'h2e5b; 14'h166a: x = 16'h2e5a; 14'h166b: x = 16'h2e59; 14'h166c: x = 16'h2e58; 14'h166d: x = 16'h2e57; 14'h166e: x = 16'h2e56; 14'h166f: x = 16'h2e55; 14'h1670: x = 16'h2e54; 14'h1671: x = 16'h2e53; 14'h1672: x = 16'h2e52; 14'h1673: x = 16'h2e51; 14'h1674: x = 16'h2e50; 14'h1675: x = 16'h2e4f; 14'h1676: x = 16'h2e4e; 14'h1677: x = 16'h2e4d; 14'h1678: x = 16'h2e4c; 14'h1679: x = 16'h2e4c; 14'h167a: x = 16'h2e4b; 14'h167b: x = 16'h2e4a; 14'h167c: x = 16'h2e49; 14'h167d: x = 16'h2e48; 14'h167e: x = 16'h2e47; 14'h167f: x = 16'h2e46; 14'h1680: x = 16'h2e45; 14'h1681: x = 16'h2e44; 14'h1682: x = 16'h2e43; 14'h1683: x = 16'h2e42; 14'h1684: x = 16'h2e41; 14'h1685: x = 16'h2e40; 14'h1686: x = 16'h2e3f; 14'h1687: x = 16'h2e3e; 14'h1688: x = 16'h2e3d; 14'h1689: x = 16'h2e3c; 14'h168a: x = 16'h2e3b; 14'h168b: x = 16'h2e3a; 14'h168c: x = 16'h2e39; 14'h168d: x = 16'h2e38; 14'h168e: x = 16'h2e37; 14'h168f: x = 16'h2e36; 14'h1690: x = 16'h2e35; 14'h1691: x = 16'h2e34; 14'h1692: x = 16'h2e33; 14'h1693: x = 16'h2e32; 14'h1694: x = 16'h2e31; 14'h1695: x = 16'h2e30; 14'h1696: x = 16'h2e2f; 14'h1697: x = 16'h2e2e; 14'h1698: x = 16'h2e2d; 14'h1699: x = 16'h2e2c; 14'h169a: x = 16'h2e2b; 14'h169b: x = 16'h2e2a; 14'h169c: x = 16'h2e29; 14'h169d: x = 16'h2e28; 14'h169e: x = 16'h2e27; 14'h169f: x = 16'h2e26; 14'h16a0: x = 16'h2e25; 14'h16a1: x = 16'h2e24; 14'h16a2: x = 16'h2e23; 14'h16a3: x = 16'h2e22; 14'h16a4: x = 16'h2e21; 14'h16a5: x = 16'h2e20; 14'h16a6: x = 16'h2e1f; 14'h16a7: x = 16'h2e1e; 14'h16a8: x = 16'h2e1d; 14'h16a9: x = 16'h2e1c; 14'h16aa: x = 16'h2e1b; 14'h16ab: x = 16'h2e1a; 14'h16ac: x = 16'h2e19; 14'h16ad: x = 16'h2e18; 14'h16ae: x = 16'h2e17; 14'h16af: x = 16'h2e16; 14'h16b0: x = 16'h2e16; 14'h16b1: x = 16'h2e15; 14'h16b2: x = 16'h2e14; 14'h16b3: x = 16'h2e13; 14'h16b4: x = 16'h2e12; 14'h16b5: x = 16'h2e11; 14'h16b6: x = 16'h2e10; 14'h16b7: x = 16'h2e0f; 14'h16b8: x = 16'h2e0e; 14'h16b9: x = 16'h2e0d; 14'h16ba: x = 16'h2e0c; 14'h16bb: x = 16'h2e0b; 14'h16bc: x = 16'h2e0a; 14'h16bd: x = 16'h2e09; 14'h16be: x = 16'h2e08; 14'h16bf: x = 16'h2e07; 14'h16c0: x = 16'h2e06; 14'h16c1: x = 16'h2e05; 14'h16c2: x = 16'h2e04; 14'h16c3: x = 16'h2e03; 14'h16c4: x = 16'h2e02; 14'h16c5: x = 16'h2e01; 14'h16c6: x = 16'h2e00; 14'h16c7: x = 16'h2dff; 14'h16c8: x = 16'h2dfe; 14'h16c9: x = 16'h2dfd; 14'h16ca: x = 16'h2dfc; 14'h16cb: x = 16'h2dfb; 14'h16cc: x = 16'h2dfa; 14'h16cd: x = 16'h2df9; 14'h16ce: x = 16'h2df8; 14'h16cf: x = 16'h2df7; 14'h16d0: x = 16'h2df6; 14'h16d1: x = 16'h2df5; 14'h16d2: x = 16'h2df4; 14'h16d3: x = 16'h2df3; 14'h16d4: x = 16'h2df2; 14'h16d5: x = 16'h2df1; 14'h16d6: x = 16'h2df0; 14'h16d7: x = 16'h2def; 14'h16d8: x = 16'h2dee; 14'h16d9: x = 16'h2ded; 14'h16da: x = 16'h2dec; 14'h16db: x = 16'h2deb; 14'h16dc: x = 16'h2deb; 14'h16dd: x = 16'h2dea; 14'h16de: x = 16'h2de9; 14'h16df: x = 16'h2de8; 14'h16e0: x = 16'h2de7; 14'h16e1: x = 16'h2de6; 14'h16e2: x = 16'h2de5; 14'h16e3: x = 16'h2de4; 14'h16e4: x = 16'h2de3; 14'h16e5: x = 16'h2de2; 14'h16e6: x = 16'h2de1; 14'h16e7: x = 16'h2de0; 14'h16e8: x = 16'h2ddf; 14'h16e9: x = 16'h2dde; 14'h16ea: x = 16'h2ddd; 14'h16eb: x = 16'h2ddc; 14'h16ec: x = 16'h2ddb; 14'h16ed: x = 16'h2dda; 14'h16ee: x = 16'h2dd9; 14'h16ef: x = 16'h2dd8; 14'h16f0: x = 16'h2dd7; 14'h16f1: x = 16'h2dd6; 14'h16f2: x = 16'h2dd5; 14'h16f3: x = 16'h2dd4; 14'h16f4: x = 16'h2dd3; 14'h16f5: x = 16'h2dd2; 14'h16f6: x = 16'h2dd1; 14'h16f7: x = 16'h2dd0; 14'h16f8: x = 16'h2dcf; 14'h16f9: x = 16'h2dce; 14'h16fa: x = 16'h2dcd; 14'h16fb: x = 16'h2dcc; 14'h16fc: x = 16'h2dcb; 14'h16fd: x = 16'h2dca; 14'h16fe: x = 16'h2dc9; 14'h16ff: x = 16'h2dc8; 14'h1700: x = 16'h2dc7; 14'h1701: x = 16'h2dc6; 14'h1702: x = 16'h2dc5; 14'h1703: x = 16'h2dc5; 14'h1704: x = 16'h2dc4; 14'h1705: x = 16'h2dc3; 14'h1706: x = 16'h2dc2; 14'h1707: x = 16'h2dc1; 14'h1708: x = 16'h2dc0; 14'h1709: x = 16'h2dbf; 14'h170a: x = 16'h2dbe; 14'h170b: x = 16'h2dbd; 14'h170c: x = 16'h2dbc; 14'h170d: x = 16'h2dbb; 14'h170e: x = 16'h2dba; 14'h170f: x = 16'h2db9; 14'h1710: x = 16'h2db8; 14'h1711: x = 16'h2db7; 14'h1712: x = 16'h2db6; 14'h1713: x = 16'h2db5; 14'h1714: x = 16'h2db4; 14'h1715: x = 16'h2db3; 14'h1716: x = 16'h2db2; 14'h1717: x = 16'h2db1; 14'h1718: x = 16'h2db0; 14'h1719: x = 16'h2daf; 14'h171a: x = 16'h2dae; 14'h171b: x = 16'h2dad; 14'h171c: x = 16'h2dac; 14'h171d: x = 16'h2dab; 14'h171e: x = 16'h2daa; 14'h171f: x = 16'h2da9; 14'h1720: x = 16'h2da8; 14'h1721: x = 16'h2da7; 14'h1722: x = 16'h2da6; 14'h1723: x = 16'h2da5; 14'h1724: x = 16'h2da4; 14'h1725: x = 16'h2da4; 14'h1726: x = 16'h2da3; 14'h1727: x = 16'h2da2; 14'h1728: x = 16'h2da1; 14'h1729: x = 16'h2da0; 14'h172a: x = 16'h2d9f; 14'h172b: x = 16'h2d9e; 14'h172c: x = 16'h2d9d; 14'h172d: x = 16'h2d9c; 14'h172e: x = 16'h2d9b; 14'h172f: x = 16'h2d9a; 14'h1730: x = 16'h2d99; 14'h1731: x = 16'h2d98; 14'h1732: x = 16'h2d97; 14'h1733: x = 16'h2d96; 14'h1734: x = 16'h2d95; 14'h1735: x = 16'h2d94; 14'h1736: x = 16'h2d93; 14'h1737: x = 16'h2d92; 14'h1738: x = 16'h2d91; 14'h1739: x = 16'h2d90; 14'h173a: x = 16'h2d8f; 14'h173b: x = 16'h2d8e; 14'h173c: x = 16'h2d8d; 14'h173d: x = 16'h2d8c; 14'h173e: x = 16'h2d8b; 14'h173f: x = 16'h2d8a; 14'h1740: x = 16'h2d89; 14'h1741: x = 16'h2d88; 14'h1742: x = 16'h2d87; 14'h1743: x = 16'h2d86; 14'h1744: x = 16'h2d86; 14'h1745: x = 16'h2d85; 14'h1746: x = 16'h2d84; 14'h1747: x = 16'h2d83; 14'h1748: x = 16'h2d82; 14'h1749: x = 16'h2d81; 14'h174a: x = 16'h2d80; 14'h174b: x = 16'h2d7f; 14'h174c: x = 16'h2d7e; 14'h174d: x = 16'h2d7d; 14'h174e: x = 16'h2d7c; 14'h174f: x = 16'h2d7b; 14'h1750: x = 16'h2d7a; 14'h1751: x = 16'h2d79; 14'h1752: x = 16'h2d78; 14'h1753: x = 16'h2d77; 14'h1754: x = 16'h2d76; 14'h1755: x = 16'h2d75; 14'h1756: x = 16'h2d74; 14'h1757: x = 16'h2d73; 14'h1758: x = 16'h2d72; 14'h1759: x = 16'h2d71; 14'h175a: x = 16'h2d70; 14'h175b: x = 16'h2d6f; 14'h175c: x = 16'h2d6e; 14'h175d: x = 16'h2d6d; 14'h175e: x = 16'h2d6c; 14'h175f: x = 16'h2d6b; 14'h1760: x = 16'h2d6a; 14'h1761: x = 16'h2d69; 14'h1762: x = 16'h2d69; 14'h1763: x = 16'h2d68; 14'h1764: x = 16'h2d67; 14'h1765: x = 16'h2d66; 14'h1766: x = 16'h2d65; 14'h1767: x = 16'h2d64; 14'h1768: x = 16'h2d63; 14'h1769: x = 16'h2d62; 14'h176a: x = 16'h2d61; 14'h176b: x = 16'h2d60; 14'h176c: x = 16'h2d5f; 14'h176d: x = 16'h2d5e; 14'h176e: x = 16'h2d5d; 14'h176f: x = 16'h2d5c; 14'h1770: x = 16'h2d5b; 14'h1771: x = 16'h2d5a; 14'h1772: x = 16'h2d59; 14'h1773: x = 16'h2d58; 14'h1774: x = 16'h2d57; 14'h1775: x = 16'h2d56; 14'h1776: x = 16'h2d55; 14'h1777: x = 16'h2d54; 14'h1778: x = 16'h2d53; 14'h1779: x = 16'h2d52; 14'h177a: x = 16'h2d51; 14'h177b: x = 16'h2d50; 14'h177c: x = 16'h2d4f; 14'h177d: x = 16'h2d4f; 14'h177e: x = 16'h2d4e; 14'h177f: x = 16'h2d4d; 14'h1780: x = 16'h2d4c; 14'h1781: x = 16'h2d4b; 14'h1782: x = 16'h2d4a; 14'h1783: x = 16'h2d49; 14'h1784: x = 16'h2d48; 14'h1785: x = 16'h2d47; 14'h1786: x = 16'h2d46; 14'h1787: x = 16'h2d45; 14'h1788: x = 16'h2d44; 14'h1789: x = 16'h2d43; 14'h178a: x = 16'h2d42; 14'h178b: x = 16'h2d41; 14'h178c: x = 16'h2d40; 14'h178d: x = 16'h2d3f; 14'h178e: x = 16'h2d3e; 14'h178f: x = 16'h2d3d; 14'h1790: x = 16'h2d3c; 14'h1791: x = 16'h2d3b; 14'h1792: x = 16'h2d3a; 14'h1793: x = 16'h2d39; 14'h1794: x = 16'h2d38; 14'h1795: x = 16'h2d37; 14'h1796: x = 16'h2d36; 14'h1797: x = 16'h2d36; 14'h1798: x = 16'h2d35; 14'h1799: x = 16'h2d34; 14'h179a: x = 16'h2d33; 14'h179b: x = 16'h2d32; 14'h179c: x = 16'h2d31; 14'h179d: x = 16'h2d30; 14'h179e: x = 16'h2d2f; 14'h179f: x = 16'h2d2e; 14'h17a0: x = 16'h2d2d; 14'h17a1: x = 16'h2d2c; 14'h17a2: x = 16'h2d2b; 14'h17a3: x = 16'h2d2a; 14'h17a4: x = 16'h2d29; 14'h17a5: x = 16'h2d28; 14'h17a6: x = 16'h2d27; 14'h17a7: x = 16'h2d26; 14'h17a8: x = 16'h2d25; 14'h17a9: x = 16'h2d24; 14'h17aa: x = 16'h2d23; 14'h17ab: x = 16'h2d22; 14'h17ac: x = 16'h2d21; 14'h17ad: x = 16'h2d20; 14'h17ae: x = 16'h2d1f; 14'h17af: x = 16'h2d1f; 14'h17b0: x = 16'h2d1e; 14'h17b1: x = 16'h2d1d; 14'h17b2: x = 16'h2d1c; 14'h17b3: x = 16'h2d1b; 14'h17b4: x = 16'h2d1a; 14'h17b5: x = 16'h2d19; 14'h17b6: x = 16'h2d18; 14'h17b7: x = 16'h2d17; 14'h17b8: x = 16'h2d16; 14'h17b9: x = 16'h2d15; 14'h17ba: x = 16'h2d14; 14'h17bb: x = 16'h2d13; 14'h17bc: x = 16'h2d12; 14'h17bd: x = 16'h2d11; 14'h17be: x = 16'h2d10; 14'h17bf: x = 16'h2d0f; 14'h17c0: x = 16'h2d0e; 14'h17c1: x = 16'h2d0d; 14'h17c2: x = 16'h2d0c; 14'h17c3: x = 16'h2d0b; 14'h17c4: x = 16'h2d0a; 14'h17c5: x = 16'h2d09; 14'h17c6: x = 16'h2d08; 14'h17c7: x = 16'h2d08; 14'h17c8: x = 16'h2d07; 14'h17c9: x = 16'h2d06; 14'h17ca: x = 16'h2d05; 14'h17cb: x = 16'h2d04; 14'h17cc: x = 16'h2d03; 14'h17cd: x = 16'h2d02; 14'h17ce: x = 16'h2d01; 14'h17cf: x = 16'h2d00; 14'h17d0: x = 16'h2cff; 14'h17d1: x = 16'h2cfe; 14'h17d2: x = 16'h2cfd; 14'h17d3: x = 16'h2cfc; 14'h17d4: x = 16'h2cfb; 14'h17d5: x = 16'h2cfa; 14'h17d6: x = 16'h2cf9; 14'h17d7: x = 16'h2cf8; 14'h17d8: x = 16'h2cf7; 14'h17d9: x = 16'h2cf6; 14'h17da: x = 16'h2cf5; 14'h17db: x = 16'h2cf4; 14'h17dc: x = 16'h2cf3; 14'h17dd: x = 16'h2cf3; 14'h17de: x = 16'h2cf2; 14'h17df: x = 16'h2cf1; 14'h17e0: x = 16'h2cf0; 14'h17e1: x = 16'h2cef; 14'h17e2: x = 16'h2cee; 14'h17e3: x = 16'h2ced; 14'h17e4: x = 16'h2cec; 14'h17e5: x = 16'h2ceb; 14'h17e6: x = 16'h2cea; 14'h17e7: x = 16'h2ce9; 14'h17e8: x = 16'h2ce8; 14'h17e9: x = 16'h2ce7; 14'h17ea: x = 16'h2ce6; 14'h17eb: x = 16'h2ce5; 14'h17ec: x = 16'h2ce4; 14'h17ed: x = 16'h2ce3; 14'h17ee: x = 16'h2ce2; 14'h17ef: x = 16'h2ce1; 14'h17f0: x = 16'h2ce0; 14'h17f1: x = 16'h2cdf; 14'h17f2: x = 16'h2cde; 14'h17f3: x = 16'h2cde; 14'h17f4: x = 16'h2cdd; 14'h17f5: x = 16'h2cdc; 14'h17f6: x = 16'h2cdb; 14'h17f7: x = 16'h2cda; 14'h17f8: x = 16'h2cd9; 14'h17f9: x = 16'h2cd8; 14'h17fa: x = 16'h2cd7; 14'h17fb: x = 16'h2cd6; 14'h17fc: x = 16'h2cd5; 14'h17fd: x = 16'h2cd4; 14'h17fe: x = 16'h2cd3; 14'h17ff: x = 16'h2cd2; 14'h1800: x = 16'h2cd1; 14'h1801: x = 16'h2cd0; 14'h1802: x = 16'h2ccf; 14'h1803: x = 16'h2cce; 14'h1804: x = 16'h2ccd; 14'h1805: x = 16'h2ccc; 14'h1806: x = 16'h2ccb; 14'h1807: x = 16'h2cca; 14'h1808: x = 16'h2cca; 14'h1809: x = 16'h2cc9; 14'h180a: x = 16'h2cc8; 14'h180b: x = 16'h2cc7; 14'h180c: x = 16'h2cc6; 14'h180d: x = 16'h2cc5; 14'h180e: x = 16'h2cc4; 14'h180f: x = 16'h2cc3; 14'h1810: x = 16'h2cc2; 14'h1811: x = 16'h2cc1; 14'h1812: x = 16'h2cc0; 14'h1813: x = 16'h2cbf; 14'h1814: x = 16'h2cbe; 14'h1815: x = 16'h2cbd; 14'h1816: x = 16'h2cbc; 14'h1817: x = 16'h2cbb; 14'h1818: x = 16'h2cba; 14'h1819: x = 16'h2cb9; 14'h181a: x = 16'h2cb8; 14'h181b: x = 16'h2cb7; 14'h181c: x = 16'h2cb7; 14'h181d: x = 16'h2cb6; 14'h181e: x = 16'h2cb5; 14'h181f: x = 16'h2cb4; 14'h1820: x = 16'h2cb3; 14'h1821: x = 16'h2cb2; 14'h1822: x = 16'h2cb1; 14'h1823: x = 16'h2cb0; 14'h1824: x = 16'h2caf; 14'h1825: x = 16'h2cae; 14'h1826: x = 16'h2cad; 14'h1827: x = 16'h2cac; 14'h1828: x = 16'h2cab; 14'h1829: x = 16'h2caa; 14'h182a: x = 16'h2ca9; 14'h182b: x = 16'h2ca8; 14'h182c: x = 16'h2ca7; 14'h182d: x = 16'h2ca6; 14'h182e: x = 16'h2ca5; 14'h182f: x = 16'h2ca4; 14'h1830: x = 16'h2ca4; 14'h1831: x = 16'h2ca3; 14'h1832: x = 16'h2ca2; 14'h1833: x = 16'h2ca1; 14'h1834: x = 16'h2ca0; 14'h1835: x = 16'h2c9f; 14'h1836: x = 16'h2c9e; 14'h1837: x = 16'h2c9d; 14'h1838: x = 16'h2c9c; 14'h1839: x = 16'h2c9b; 14'h183a: x = 16'h2c9a; 14'h183b: x = 16'h2c99; 14'h183c: x = 16'h2c98; 14'h183d: x = 16'h2c97; 14'h183e: x = 16'h2c96; 14'h183f: x = 16'h2c95; 14'h1840: x = 16'h2c94; 14'h1841: x = 16'h2c93; 14'h1842: x = 16'h2c92; 14'h1843: x = 16'h2c92; 14'h1844: x = 16'h2c91; 14'h1845: x = 16'h2c90; 14'h1846: x = 16'h2c8f; 14'h1847: x = 16'h2c8e; 14'h1848: x = 16'h2c8d; 14'h1849: x = 16'h2c8c; 14'h184a: x = 16'h2c8b; 14'h184b: x = 16'h2c8a; 14'h184c: x = 16'h2c89; 14'h184d: x = 16'h2c88; 14'h184e: x = 16'h2c87; 14'h184f: x = 16'h2c86; 14'h1850: x = 16'h2c85; 14'h1851: x = 16'h2c84; 14'h1852: x = 16'h2c83; 14'h1853: x = 16'h2c82; 14'h1854: x = 16'h2c81; 14'h1855: x = 16'h2c81; 14'h1856: x = 16'h2c80; 14'h1857: x = 16'h2c7f; 14'h1858: x = 16'h2c7e; 14'h1859: x = 16'h2c7d; 14'h185a: x = 16'h2c7c; 14'h185b: x = 16'h2c7b; 14'h185c: x = 16'h2c7a; 14'h185d: x = 16'h2c79; 14'h185e: x = 16'h2c78; 14'h185f: x = 16'h2c77; 14'h1860: x = 16'h2c76; 14'h1861: x = 16'h2c75; 14'h1862: x = 16'h2c74; 14'h1863: x = 16'h2c73; 14'h1864: x = 16'h2c72; 14'h1865: x = 16'h2c71; 14'h1866: x = 16'h2c70; 14'h1867: x = 16'h2c6f; 14'h1868: x = 16'h2c6f; 14'h1869: x = 16'h2c6e; 14'h186a: x = 16'h2c6d; 14'h186b: x = 16'h2c6c; 14'h186c: x = 16'h2c6b; 14'h186d: x = 16'h2c6a; 14'h186e: x = 16'h2c69; 14'h186f: x = 16'h2c68; 14'h1870: x = 16'h2c67; 14'h1871: x = 16'h2c66; 14'h1872: x = 16'h2c65; 14'h1873: x = 16'h2c64; 14'h1874: x = 16'h2c63; 14'h1875: x = 16'h2c62; 14'h1876: x = 16'h2c61; 14'h1877: x = 16'h2c60; 14'h1878: x = 16'h2c5f; 14'h1879: x = 16'h2c5f; 14'h187a: x = 16'h2c5e; 14'h187b: x = 16'h2c5d; 14'h187c: x = 16'h2c5c; 14'h187d: x = 16'h2c5b; 14'h187e: x = 16'h2c5a; 14'h187f: x = 16'h2c59; 14'h1880: x = 16'h2c58; 14'h1881: x = 16'h2c57; 14'h1882: x = 16'h2c56; 14'h1883: x = 16'h2c55; 14'h1884: x = 16'h2c54; 14'h1885: x = 16'h2c53; 14'h1886: x = 16'h2c52; 14'h1887: x = 16'h2c51; 14'h1888: x = 16'h2c50; 14'h1889: x = 16'h2c4f; 14'h188a: x = 16'h2c4e; 14'h188b: x = 16'h2c4e; 14'h188c: x = 16'h2c4d; 14'h188d: x = 16'h2c4c; 14'h188e: x = 16'h2c4b; 14'h188f: x = 16'h2c4a; 14'h1890: x = 16'h2c49; 14'h1891: x = 16'h2c48; 14'h1892: x = 16'h2c47; 14'h1893: x = 16'h2c46; 14'h1894: x = 16'h2c45; 14'h1895: x = 16'h2c44; 14'h1896: x = 16'h2c43; 14'h1897: x = 16'h2c42; 14'h1898: x = 16'h2c41; 14'h1899: x = 16'h2c40; 14'h189a: x = 16'h2c3f; 14'h189b: x = 16'h2c3e; 14'h189c: x = 16'h2c3e; 14'h189d: x = 16'h2c3d; 14'h189e: x = 16'h2c3c; 14'h189f: x = 16'h2c3b; 14'h18a0: x = 16'h2c3a; 14'h18a1: x = 16'h2c39; 14'h18a2: x = 16'h2c38; 14'h18a3: x = 16'h2c37; 14'h18a4: x = 16'h2c36; 14'h18a5: x = 16'h2c35; 14'h18a6: x = 16'h2c34; 14'h18a7: x = 16'h2c33; 14'h18a8: x = 16'h2c32; 14'h18a9: x = 16'h2c31; 14'h18aa: x = 16'h2c30; 14'h18ab: x = 16'h2c2f; 14'h18ac: x = 16'h2c2f; 14'h18ad: x = 16'h2c2e; 14'h18ae: x = 16'h2c2d; 14'h18af: x = 16'h2c2c; 14'h18b0: x = 16'h2c2b; 14'h18b1: x = 16'h2c2a; 14'h18b2: x = 16'h2c29; 14'h18b3: x = 16'h2c28; 14'h18b4: x = 16'h2c27; 14'h18b5: x = 16'h2c26; 14'h18b6: x = 16'h2c25; 14'h18b7: x = 16'h2c24; 14'h18b8: x = 16'h2c23; 14'h18b9: x = 16'h2c22; 14'h18ba: x = 16'h2c21; 14'h18bb: x = 16'h2c20; 14'h18bc: x = 16'h2c1f; 14'h18bd: x = 16'h2c1f; 14'h18be: x = 16'h2c1e; 14'h18bf: x = 16'h2c1d; 14'h18c0: x = 16'h2c1c; 14'h18c1: x = 16'h2c1b; 14'h18c2: x = 16'h2c1a; 14'h18c3: x = 16'h2c19; 14'h18c4: x = 16'h2c18; 14'h18c5: x = 16'h2c17; 14'h18c6: x = 16'h2c16; 14'h18c7: x = 16'h2c15; 14'h18c8: x = 16'h2c14; 14'h18c9: x = 16'h2c13; 14'h18ca: x = 16'h2c12; 14'h18cb: x = 16'h2c11; 14'h18cc: x = 16'h2c10; 14'h18cd: x = 16'h2c10; 14'h18ce: x = 16'h2c0f; 14'h18cf: x = 16'h2c0e; 14'h18d0: x = 16'h2c0d; 14'h18d1: x = 16'h2c0c; 14'h18d2: x = 16'h2c0b; 14'h18d3: x = 16'h2c0a; 14'h18d4: x = 16'h2c09; 14'h18d5: x = 16'h2c08; 14'h18d6: x = 16'h2c07; 14'h18d7: x = 16'h2c06; 14'h18d8: x = 16'h2c05; 14'h18d9: x = 16'h2c04; 14'h18da: x = 16'h2c03; 14'h18db: x = 16'h2c02; 14'h18dc: x = 16'h2c01; 14'h18dd: x = 16'h2c01; 14'h18de: x = 16'h2c00; 14'h18df: x = 16'h2bff; 14'h18e0: x = 16'h2bfe; 14'h18e1: x = 16'h2bfd; 14'h18e2: x = 16'h2bfc; 14'h18e3: x = 16'h2bfb; 14'h18e4: x = 16'h2bfa; 14'h18e5: x = 16'h2bf9; 14'h18e6: x = 16'h2bf8; 14'h18e7: x = 16'h2bf7; 14'h18e8: x = 16'h2bf6; 14'h18e9: x = 16'h2bf5; 14'h18ea: x = 16'h2bf4; 14'h18eb: x = 16'h2bf3; 14'h18ec: x = 16'h2bf3; 14'h18ed: x = 16'h2bf2; 14'h18ee: x = 16'h2bf1; 14'h18ef: x = 16'h2bf0; 14'h18f0: x = 16'h2bef; 14'h18f1: x = 16'h2bee; 14'h18f2: x = 16'h2bed; 14'h18f3: x = 16'h2bec; 14'h18f4: x = 16'h2beb; 14'h18f5: x = 16'h2bea; 14'h18f6: x = 16'h2be9; 14'h18f7: x = 16'h2be8; 14'h18f8: x = 16'h2be7; 14'h18f9: x = 16'h2be6; 14'h18fa: x = 16'h2be5; 14'h18fb: x = 16'h2be5; 14'h18fc: x = 16'h2be4; 14'h18fd: x = 16'h2be3; 14'h18fe: x = 16'h2be2; 14'h18ff: x = 16'h2be1; 14'h1900: x = 16'h2be0; 14'h1901: x = 16'h2bdf; 14'h1902: x = 16'h2bde; 14'h1903: x = 16'h2bdd; 14'h1904: x = 16'h2bdc; 14'h1905: x = 16'h2bdb; 14'h1906: x = 16'h2bda; 14'h1907: x = 16'h2bd9; 14'h1908: x = 16'h2bd8; 14'h1909: x = 16'h2bd7; 14'h190a: x = 16'h2bd7; 14'h190b: x = 16'h2bd6; 14'h190c: x = 16'h2bd5; 14'h190d: x = 16'h2bd4; 14'h190e: x = 16'h2bd3; 14'h190f: x = 16'h2bd2; 14'h1910: x = 16'h2bd1; 14'h1911: x = 16'h2bd0; 14'h1912: x = 16'h2bcf; 14'h1913: x = 16'h2bce; 14'h1914: x = 16'h2bcd; 14'h1915: x = 16'h2bcc; 14'h1916: x = 16'h2bcb; 14'h1917: x = 16'h2bca; 14'h1918: x = 16'h2bc9; 14'h1919: x = 16'h2bc9; 14'h191a: x = 16'h2bc8; 14'h191b: x = 16'h2bc7; 14'h191c: x = 16'h2bc6; 14'h191d: x = 16'h2bc5; 14'h191e: x = 16'h2bc4; 14'h191f: x = 16'h2bc3; 14'h1920: x = 16'h2bc2; 14'h1921: x = 16'h2bc1; 14'h1922: x = 16'h2bc0; 14'h1923: x = 16'h2bbf; 14'h1924: x = 16'h2bbe; 14'h1925: x = 16'h2bbd; 14'h1926: x = 16'h2bbc; 14'h1927: x = 16'h2bbb; 14'h1928: x = 16'h2bbb; 14'h1929: x = 16'h2bba; 14'h192a: x = 16'h2bb9; 14'h192b: x = 16'h2bb8; 14'h192c: x = 16'h2bb7; 14'h192d: x = 16'h2bb6; 14'h192e: x = 16'h2bb5; 14'h192f: x = 16'h2bb4; 14'h1930: x = 16'h2bb3; 14'h1931: x = 16'h2bb2; 14'h1932: x = 16'h2bb1; 14'h1933: x = 16'h2bb0; 14'h1934: x = 16'h2baf; 14'h1935: x = 16'h2bae; 14'h1936: x = 16'h2bae; 14'h1937: x = 16'h2bad; 14'h1938: x = 16'h2bac; 14'h1939: x = 16'h2bab; 14'h193a: x = 16'h2baa; 14'h193b: x = 16'h2ba9; 14'h193c: x = 16'h2ba8; 14'h193d: x = 16'h2ba7; 14'h193e: x = 16'h2ba6; 14'h193f: x = 16'h2ba5; 14'h1940: x = 16'h2ba4; 14'h1941: x = 16'h2ba3; 14'h1942: x = 16'h2ba2; 14'h1943: x = 16'h2ba1; 14'h1944: x = 16'h2ba1; 14'h1945: x = 16'h2ba0; 14'h1946: x = 16'h2b9f; 14'h1947: x = 16'h2b9e; 14'h1948: x = 16'h2b9d; 14'h1949: x = 16'h2b9c; 14'h194a: x = 16'h2b9b; 14'h194b: x = 16'h2b9a; 14'h194c: x = 16'h2b99; 14'h194d: x = 16'h2b98; 14'h194e: x = 16'h2b97; 14'h194f: x = 16'h2b96; 14'h1950: x = 16'h2b95; 14'h1951: x = 16'h2b94; 14'h1952: x = 16'h2b94; 14'h1953: x = 16'h2b93; 14'h1954: x = 16'h2b92; 14'h1955: x = 16'h2b91; 14'h1956: x = 16'h2b90; 14'h1957: x = 16'h2b8f; 14'h1958: x = 16'h2b8e; 14'h1959: x = 16'h2b8d; 14'h195a: x = 16'h2b8c; 14'h195b: x = 16'h2b8b; 14'h195c: x = 16'h2b8a; 14'h195d: x = 16'h2b89; 14'h195e: x = 16'h2b88; 14'h195f: x = 16'h2b87; 14'h1960: x = 16'h2b87; 14'h1961: x = 16'h2b86; 14'h1962: x = 16'h2b85; 14'h1963: x = 16'h2b84; 14'h1964: x = 16'h2b83; 14'h1965: x = 16'h2b82; 14'h1966: x = 16'h2b81; 14'h1967: x = 16'h2b80; 14'h1968: x = 16'h2b7f; 14'h1969: x = 16'h2b7e; 14'h196a: x = 16'h2b7d; 14'h196b: x = 16'h2b7c; 14'h196c: x = 16'h2b7b; 14'h196d: x = 16'h2b7a; 14'h196e: x = 16'h2b7a; 14'h196f: x = 16'h2b79; 14'h1970: x = 16'h2b78; 14'h1971: x = 16'h2b77; 14'h1972: x = 16'h2b76; 14'h1973: x = 16'h2b75; 14'h1974: x = 16'h2b74; 14'h1975: x = 16'h2b73; 14'h1976: x = 16'h2b72; 14'h1977: x = 16'h2b71; 14'h1978: x = 16'h2b70; 14'h1979: x = 16'h2b6f; 14'h197a: x = 16'h2b6e; 14'h197b: x = 16'h2b6e; 14'h197c: x = 16'h2b6d; 14'h197d: x = 16'h2b6c; 14'h197e: x = 16'h2b6b; 14'h197f: x = 16'h2b6a; 14'h1980: x = 16'h2b69; 14'h1981: x = 16'h2b68; 14'h1982: x = 16'h2b67; 14'h1983: x = 16'h2b66; 14'h1984: x = 16'h2b65; 14'h1985: x = 16'h2b64; 14'h1986: x = 16'h2b63; 14'h1987: x = 16'h2b62; 14'h1988: x = 16'h2b62; 14'h1989: x = 16'h2b61; 14'h198a: x = 16'h2b60; 14'h198b: x = 16'h2b5f; 14'h198c: x = 16'h2b5e; 14'h198d: x = 16'h2b5d; 14'h198e: x = 16'h2b5c; 14'h198f: x = 16'h2b5b; 14'h1990: x = 16'h2b5a; 14'h1991: x = 16'h2b59; 14'h1992: x = 16'h2b58; 14'h1993: x = 16'h2b57; 14'h1994: x = 16'h2b56; 14'h1995: x = 16'h2b55; 14'h1996: x = 16'h2b55; 14'h1997: x = 16'h2b54; 14'h1998: x = 16'h2b53; 14'h1999: x = 16'h2b52; 14'h199a: x = 16'h2b51; 14'h199b: x = 16'h2b50; 14'h199c: x = 16'h2b4f; 14'h199d: x = 16'h2b4e; 14'h199e: x = 16'h2b4d; 14'h199f: x = 16'h2b4c; 14'h19a0: x = 16'h2b4b; 14'h19a1: x = 16'h2b4a; 14'h19a2: x = 16'h2b49; 14'h19a3: x = 16'h2b49; 14'h19a4: x = 16'h2b48; 14'h19a5: x = 16'h2b47; 14'h19a6: x = 16'h2b46; 14'h19a7: x = 16'h2b45; 14'h19a8: x = 16'h2b44; 14'h19a9: x = 16'h2b43; 14'h19aa: x = 16'h2b42; 14'h19ab: x = 16'h2b41; 14'h19ac: x = 16'h2b40; 14'h19ad: x = 16'h2b3f; 14'h19ae: x = 16'h2b3e; 14'h19af: x = 16'h2b3e; 14'h19b0: x = 16'h2b3d; 14'h19b1: x = 16'h2b3c; 14'h19b2: x = 16'h2b3b; 14'h19b3: x = 16'h2b3a; 14'h19b4: x = 16'h2b39; 14'h19b5: x = 16'h2b38; 14'h19b6: x = 16'h2b37; 14'h19b7: x = 16'h2b36; 14'h19b8: x = 16'h2b35; 14'h19b9: x = 16'h2b34; 14'h19ba: x = 16'h2b33; 14'h19bb: x = 16'h2b32; 14'h19bc: x = 16'h2b32; 14'h19bd: x = 16'h2b31; 14'h19be: x = 16'h2b30; 14'h19bf: x = 16'h2b2f; 14'h19c0: x = 16'h2b2e; 14'h19c1: x = 16'h2b2d; 14'h19c2: x = 16'h2b2c; 14'h19c3: x = 16'h2b2b; 14'h19c4: x = 16'h2b2a; 14'h19c5: x = 16'h2b29; 14'h19c6: x = 16'h2b28; 14'h19c7: x = 16'h2b27; 14'h19c8: x = 16'h2b26; 14'h19c9: x = 16'h2b26; 14'h19ca: x = 16'h2b25; 14'h19cb: x = 16'h2b24; 14'h19cc: x = 16'h2b23; 14'h19cd: x = 16'h2b22; 14'h19ce: x = 16'h2b21; 14'h19cf: x = 16'h2b20; 14'h19d0: x = 16'h2b1f; 14'h19d1: x = 16'h2b1e; 14'h19d2: x = 16'h2b1d; 14'h19d3: x = 16'h2b1c; 14'h19d4: x = 16'h2b1b; 14'h19d5: x = 16'h2b1b; 14'h19d6: x = 16'h2b1a; 14'h19d7: x = 16'h2b19; 14'h19d8: x = 16'h2b18; 14'h19d9: x = 16'h2b17; 14'h19da: x = 16'h2b16; 14'h19db: x = 16'h2b15; 14'h19dc: x = 16'h2b14; 14'h19dd: x = 16'h2b13; 14'h19de: x = 16'h2b12; 14'h19df: x = 16'h2b11; 14'h19e0: x = 16'h2b10; 14'h19e1: x = 16'h2b0f; 14'h19e2: x = 16'h2b0f; 14'h19e3: x = 16'h2b0e; 14'h19e4: x = 16'h2b0d; 14'h19e5: x = 16'h2b0c; 14'h19e6: x = 16'h2b0b; 14'h19e7: x = 16'h2b0a; 14'h19e8: x = 16'h2b09; 14'h19e9: x = 16'h2b08; 14'h19ea: x = 16'h2b07; 14'h19eb: x = 16'h2b06; 14'h19ec: x = 16'h2b05; 14'h19ed: x = 16'h2b04; 14'h19ee: x = 16'h2b04; 14'h19ef: x = 16'h2b03; 14'h19f0: x = 16'h2b02; 14'h19f1: x = 16'h2b01; 14'h19f2: x = 16'h2b00; 14'h19f3: x = 16'h2aff; 14'h19f4: x = 16'h2afe; 14'h19f5: x = 16'h2afd; 14'h19f6: x = 16'h2afc; 14'h19f7: x = 16'h2afb; 14'h19f8: x = 16'h2afa; 14'h19f9: x = 16'h2af9; 14'h19fa: x = 16'h2af9; 14'h19fb: x = 16'h2af8; 14'h19fc: x = 16'h2af7; 14'h19fd: x = 16'h2af6; 14'h19fe: x = 16'h2af5; 14'h19ff: x = 16'h2af4; 14'h1a00: x = 16'h2af3; 14'h1a01: x = 16'h2af2; 14'h1a02: x = 16'h2af1; 14'h1a03: x = 16'h2af0; 14'h1a04: x = 16'h2aef; 14'h1a05: x = 16'h2aee; 14'h1a06: x = 16'h2aee; 14'h1a07: x = 16'h2aed; 14'h1a08: x = 16'h2aec; 14'h1a09: x = 16'h2aeb; 14'h1a0a: x = 16'h2aea; 14'h1a0b: x = 16'h2ae9; 14'h1a0c: x = 16'h2ae8; 14'h1a0d: x = 16'h2ae7; 14'h1a0e: x = 16'h2ae6; 14'h1a0f: x = 16'h2ae5; 14'h1a10: x = 16'h2ae4; 14'h1a11: x = 16'h2ae3; 14'h1a12: x = 16'h2ae3; 14'h1a13: x = 16'h2ae2; 14'h1a14: x = 16'h2ae1; 14'h1a15: x = 16'h2ae0; 14'h1a16: x = 16'h2adf; 14'h1a17: x = 16'h2ade; 14'h1a18: x = 16'h2add; 14'h1a19: x = 16'h2adc; 14'h1a1a: x = 16'h2adb; 14'h1a1b: x = 16'h2ada; 14'h1a1c: x = 16'h2ad9; 14'h1a1d: x = 16'h2ad8; 14'h1a1e: x = 16'h2ad8; 14'h1a1f: x = 16'h2ad7; 14'h1a20: x = 16'h2ad6; 14'h1a21: x = 16'h2ad5; 14'h1a22: x = 16'h2ad4; 14'h1a23: x = 16'h2ad3; 14'h1a24: x = 16'h2ad2; 14'h1a25: x = 16'h2ad1; 14'h1a26: x = 16'h2ad0; 14'h1a27: x = 16'h2acf; 14'h1a28: x = 16'h2ace; 14'h1a29: x = 16'h2acd; 14'h1a2a: x = 16'h2acd; 14'h1a2b: x = 16'h2acc; 14'h1a2c: x = 16'h2acb; 14'h1a2d: x = 16'h2aca; 14'h1a2e: x = 16'h2ac9; 14'h1a2f: x = 16'h2ac8; 14'h1a30: x = 16'h2ac7; 14'h1a31: x = 16'h2ac6; 14'h1a32: x = 16'h2ac5; 14'h1a33: x = 16'h2ac4; 14'h1a34: x = 16'h2ac3; 14'h1a35: x = 16'h2ac3; 14'h1a36: x = 16'h2ac2; 14'h1a37: x = 16'h2ac1; 14'h1a38: x = 16'h2ac0; 14'h1a39: x = 16'h2abf; 14'h1a3a: x = 16'h2abe; 14'h1a3b: x = 16'h2abd; 14'h1a3c: x = 16'h2abc; 14'h1a3d: x = 16'h2abb; 14'h1a3e: x = 16'h2aba; 14'h1a3f: x = 16'h2ab9; 14'h1a40: x = 16'h2ab8; 14'h1a41: x = 16'h2ab8; 14'h1a42: x = 16'h2ab7; 14'h1a43: x = 16'h2ab6; 14'h1a44: x = 16'h2ab5; 14'h1a45: x = 16'h2ab4; 14'h1a46: x = 16'h2ab3; 14'h1a47: x = 16'h2ab2; 14'h1a48: x = 16'h2ab1; 14'h1a49: x = 16'h2ab0; 14'h1a4a: x = 16'h2aaf; 14'h1a4b: x = 16'h2aae; 14'h1a4c: x = 16'h2aae; 14'h1a4d: x = 16'h2aad; 14'h1a4e: x = 16'h2aac; 14'h1a4f: x = 16'h2aab; 14'h1a50: x = 16'h2aaa; 14'h1a51: x = 16'h2aa9; 14'h1a52: x = 16'h2aa8; 14'h1a53: x = 16'h2aa7; 14'h1a54: x = 16'h2aa6; 14'h1a55: x = 16'h2aa5; 14'h1a56: x = 16'h2aa4; 14'h1a57: x = 16'h2aa3; 14'h1a58: x = 16'h2aa3; 14'h1a59: x = 16'h2aa2; 14'h1a5a: x = 16'h2aa1; 14'h1a5b: x = 16'h2aa0; 14'h1a5c: x = 16'h2a9f; 14'h1a5d: x = 16'h2a9e; 14'h1a5e: x = 16'h2a9d; 14'h1a5f: x = 16'h2a9c; 14'h1a60: x = 16'h2a9b; 14'h1a61: x = 16'h2a9a; 14'h1a62: x = 16'h2a99; 14'h1a63: x = 16'h2a99; 14'h1a64: x = 16'h2a98; 14'h1a65: x = 16'h2a97; 14'h1a66: x = 16'h2a96; 14'h1a67: x = 16'h2a95; 14'h1a68: x = 16'h2a94; 14'h1a69: x = 16'h2a93; 14'h1a6a: x = 16'h2a92; 14'h1a6b: x = 16'h2a91; 14'h1a6c: x = 16'h2a90; 14'h1a6d: x = 16'h2a8f; 14'h1a6e: x = 16'h2a8f; 14'h1a6f: x = 16'h2a8e; 14'h1a70: x = 16'h2a8d; 14'h1a71: x = 16'h2a8c; 14'h1a72: x = 16'h2a8b; 14'h1a73: x = 16'h2a8a; 14'h1a74: x = 16'h2a89; 14'h1a75: x = 16'h2a88; 14'h1a76: x = 16'h2a87; 14'h1a77: x = 16'h2a86; 14'h1a78: x = 16'h2a85; 14'h1a79: x = 16'h2a85; 14'h1a7a: x = 16'h2a84; 14'h1a7b: x = 16'h2a83; 14'h1a7c: x = 16'h2a82; 14'h1a7d: x = 16'h2a81; 14'h1a7e: x = 16'h2a80; 14'h1a7f: x = 16'h2a7f; 14'h1a80: x = 16'h2a7e; 14'h1a81: x = 16'h2a7d; 14'h1a82: x = 16'h2a7c; 14'h1a83: x = 16'h2a7b; 14'h1a84: x = 16'h2a7b; 14'h1a85: x = 16'h2a7a; 14'h1a86: x = 16'h2a79; 14'h1a87: x = 16'h2a78; 14'h1a88: x = 16'h2a77; 14'h1a89: x = 16'h2a76; 14'h1a8a: x = 16'h2a75; 14'h1a8b: x = 16'h2a74; 14'h1a8c: x = 16'h2a73; 14'h1a8d: x = 16'h2a72; 14'h1a8e: x = 16'h2a71; 14'h1a8f: x = 16'h2a71; 14'h1a90: x = 16'h2a70; 14'h1a91: x = 16'h2a6f; 14'h1a92: x = 16'h2a6e; 14'h1a93: x = 16'h2a6d; 14'h1a94: x = 16'h2a6c; 14'h1a95: x = 16'h2a6b; 14'h1a96: x = 16'h2a6a; 14'h1a97: x = 16'h2a69; 14'h1a98: x = 16'h2a68; 14'h1a99: x = 16'h2a67; 14'h1a9a: x = 16'h2a67; 14'h1a9b: x = 16'h2a66; 14'h1a9c: x = 16'h2a65; 14'h1a9d: x = 16'h2a64; 14'h1a9e: x = 16'h2a63; 14'h1a9f: x = 16'h2a62; 14'h1aa0: x = 16'h2a61; 14'h1aa1: x = 16'h2a60; 14'h1aa2: x = 16'h2a5f; 14'h1aa3: x = 16'h2a5e; 14'h1aa4: x = 16'h2a5d; 14'h1aa5: x = 16'h2a5d; 14'h1aa6: x = 16'h2a5c; 14'h1aa7: x = 16'h2a5b; 14'h1aa8: x = 16'h2a5a; 14'h1aa9: x = 16'h2a59; 14'h1aaa: x = 16'h2a58; 14'h1aab: x = 16'h2a57; 14'h1aac: x = 16'h2a56; 14'h1aad: x = 16'h2a55; 14'h1aae: x = 16'h2a54; 14'h1aaf: x = 16'h2a53; 14'h1ab0: x = 16'h2a53; 14'h1ab1: x = 16'h2a52; 14'h1ab2: x = 16'h2a51; 14'h1ab3: x = 16'h2a50; 14'h1ab4: x = 16'h2a4f; 14'h1ab5: x = 16'h2a4e; 14'h1ab6: x = 16'h2a4d; 14'h1ab7: x = 16'h2a4c; 14'h1ab8: x = 16'h2a4b; 14'h1ab9: x = 16'h2a4a; 14'h1aba: x = 16'h2a4a; 14'h1abb: x = 16'h2a49; 14'h1abc: x = 16'h2a48; 14'h1abd: x = 16'h2a47; 14'h1abe: x = 16'h2a46; 14'h1abf: x = 16'h2a45; 14'h1ac0: x = 16'h2a44; 14'h1ac1: x = 16'h2a43; 14'h1ac2: x = 16'h2a42; 14'h1ac3: x = 16'h2a41; 14'h1ac4: x = 16'h2a40; 14'h1ac5: x = 16'h2a40; 14'h1ac6: x = 16'h2a3f; 14'h1ac7: x = 16'h2a3e; 14'h1ac8: x = 16'h2a3d; 14'h1ac9: x = 16'h2a3c; 14'h1aca: x = 16'h2a3b; 14'h1acb: x = 16'h2a3a; 14'h1acc: x = 16'h2a39; 14'h1acd: x = 16'h2a38; 14'h1ace: x = 16'h2a37; 14'h1acf: x = 16'h2a36; 14'h1ad0: x = 16'h2a36; 14'h1ad1: x = 16'h2a35; 14'h1ad2: x = 16'h2a34; 14'h1ad3: x = 16'h2a33; 14'h1ad4: x = 16'h2a32; 14'h1ad5: x = 16'h2a31; 14'h1ad6: x = 16'h2a30; 14'h1ad7: x = 16'h2a2f; 14'h1ad8: x = 16'h2a2e; 14'h1ad9: x = 16'h2a2d; 14'h1ada: x = 16'h2a2d; 14'h1adb: x = 16'h2a2c; 14'h1adc: x = 16'h2a2b; 14'h1add: x = 16'h2a2a; 14'h1ade: x = 16'h2a29; 14'h1adf: x = 16'h2a28; 14'h1ae0: x = 16'h2a27; 14'h1ae1: x = 16'h2a26; 14'h1ae2: x = 16'h2a25; 14'h1ae3: x = 16'h2a24; 14'h1ae4: x = 16'h2a23; 14'h1ae5: x = 16'h2a23; 14'h1ae6: x = 16'h2a22; 14'h1ae7: x = 16'h2a21; 14'h1ae8: x = 16'h2a20; 14'h1ae9: x = 16'h2a1f; 14'h1aea: x = 16'h2a1e; 14'h1aeb: x = 16'h2a1d; 14'h1aec: x = 16'h2a1c; 14'h1aed: x = 16'h2a1b; 14'h1aee: x = 16'h2a1a; 14'h1aef: x = 16'h2a1a; 14'h1af0: x = 16'h2a19; 14'h1af1: x = 16'h2a18; 14'h1af2: x = 16'h2a17; 14'h1af3: x = 16'h2a16; 14'h1af4: x = 16'h2a15; 14'h1af5: x = 16'h2a14; 14'h1af6: x = 16'h2a13; 14'h1af7: x = 16'h2a12; 14'h1af8: x = 16'h2a11; 14'h1af9: x = 16'h2a11; 14'h1afa: x = 16'h2a10; 14'h1afb: x = 16'h2a0f; 14'h1afc: x = 16'h2a0e; 14'h1afd: x = 16'h2a0d; 14'h1afe: x = 16'h2a0c; 14'h1aff: x = 16'h2a0b; 14'h1b00: x = 16'h2a0a; 14'h1b01: x = 16'h2a09; 14'h1b02: x = 16'h2a08; 14'h1b03: x = 16'h2a08; 14'h1b04: x = 16'h2a07; 14'h1b05: x = 16'h2a06; 14'h1b06: x = 16'h2a05; 14'h1b07: x = 16'h2a04; 14'h1b08: x = 16'h2a03; 14'h1b09: x = 16'h2a02; 14'h1b0a: x = 16'h2a01; 14'h1b0b: x = 16'h2a00; 14'h1b0c: x = 16'h29ff; 14'h1b0d: x = 16'h29fe; 14'h1b0e: x = 16'h29fe; 14'h1b0f: x = 16'h29fd; 14'h1b10: x = 16'h29fc; 14'h1b11: x = 16'h29fb; 14'h1b12: x = 16'h29fa; 14'h1b13: x = 16'h29f9; 14'h1b14: x = 16'h29f8; 14'h1b15: x = 16'h29f7; 14'h1b16: x = 16'h29f6; 14'h1b17: x = 16'h29f5; 14'h1b18: x = 16'h29f5; 14'h1b19: x = 16'h29f4; 14'h1b1a: x = 16'h29f3; 14'h1b1b: x = 16'h29f2; 14'h1b1c: x = 16'h29f1; 14'h1b1d: x = 16'h29f0; 14'h1b1e: x = 16'h29ef; 14'h1b1f: x = 16'h29ee; 14'h1b20: x = 16'h29ed; 14'h1b21: x = 16'h29ec; 14'h1b22: x = 16'h29ec; 14'h1b23: x = 16'h29eb; 14'h1b24: x = 16'h29ea; 14'h1b25: x = 16'h29e9; 14'h1b26: x = 16'h29e8; 14'h1b27: x = 16'h29e7; 14'h1b28: x = 16'h29e6; 14'h1b29: x = 16'h29e5; 14'h1b2a: x = 16'h29e4; 14'h1b2b: x = 16'h29e3; 14'h1b2c: x = 16'h29e3; 14'h1b2d: x = 16'h29e2; 14'h1b2e: x = 16'h29e1; 14'h1b2f: x = 16'h29e0; 14'h1b30: x = 16'h29df; 14'h1b31: x = 16'h29de; 14'h1b32: x = 16'h29dd; 14'h1b33: x = 16'h29dc; 14'h1b34: x = 16'h29db; 14'h1b35: x = 16'h29da; 14'h1b36: x = 16'h29da; 14'h1b37: x = 16'h29d9; 14'h1b38: x = 16'h29d8; 14'h1b39: x = 16'h29d7; 14'h1b3a: x = 16'h29d6; 14'h1b3b: x = 16'h29d5; 14'h1b3c: x = 16'h29d4; 14'h1b3d: x = 16'h29d3; 14'h1b3e: x = 16'h29d2; 14'h1b3f: x = 16'h29d1; 14'h1b40: x = 16'h29d1; 14'h1b41: x = 16'h29d0; 14'h1b42: x = 16'h29cf; 14'h1b43: x = 16'h29ce; 14'h1b44: x = 16'h29cd; 14'h1b45: x = 16'h29cc; 14'h1b46: x = 16'h29cb; 14'h1b47: x = 16'h29ca; 14'h1b48: x = 16'h29c9; 14'h1b49: x = 16'h29c9; 14'h1b4a: x = 16'h29c8; 14'h1b4b: x = 16'h29c7; 14'h1b4c: x = 16'h29c6; 14'h1b4d: x = 16'h29c5; 14'h1b4e: x = 16'h29c4; 14'h1b4f: x = 16'h29c3; 14'h1b50: x = 16'h29c2; 14'h1b51: x = 16'h29c1; 14'h1b52: x = 16'h29c0; 14'h1b53: x = 16'h29c0; 14'h1b54: x = 16'h29bf; 14'h1b55: x = 16'h29be; 14'h1b56: x = 16'h29bd; 14'h1b57: x = 16'h29bc; 14'h1b58: x = 16'h29bb; 14'h1b59: x = 16'h29ba; 14'h1b5a: x = 16'h29b9; 14'h1b5b: x = 16'h29b8; 14'h1b5c: x = 16'h29b7; 14'h1b5d: x = 16'h29b7; 14'h1b5e: x = 16'h29b6; 14'h1b5f: x = 16'h29b5; 14'h1b60: x = 16'h29b4; 14'h1b61: x = 16'h29b3; 14'h1b62: x = 16'h29b2; 14'h1b63: x = 16'h29b1; 14'h1b64: x = 16'h29b0; 14'h1b65: x = 16'h29af; 14'h1b66: x = 16'h29ae; 14'h1b67: x = 16'h29ae; 14'h1b68: x = 16'h29ad; 14'h1b69: x = 16'h29ac; 14'h1b6a: x = 16'h29ab; 14'h1b6b: x = 16'h29aa; 14'h1b6c: x = 16'h29a9; 14'h1b6d: x = 16'h29a8; 14'h1b6e: x = 16'h29a7; 14'h1b6f: x = 16'h29a6; 14'h1b70: x = 16'h29a6; 14'h1b71: x = 16'h29a5; 14'h1b72: x = 16'h29a4; 14'h1b73: x = 16'h29a3; 14'h1b74: x = 16'h29a2; 14'h1b75: x = 16'h29a1; 14'h1b76: x = 16'h29a0; 14'h1b77: x = 16'h299f; 14'h1b78: x = 16'h299e; 14'h1b79: x = 16'h299d; 14'h1b7a: x = 16'h299d; 14'h1b7b: x = 16'h299c; 14'h1b7c: x = 16'h299b; 14'h1b7d: x = 16'h299a; 14'h1b7e: x = 16'h2999; 14'h1b7f: x = 16'h2998; 14'h1b80: x = 16'h2997; 14'h1b81: x = 16'h2996; 14'h1b82: x = 16'h2995; 14'h1b83: x = 16'h2995; 14'h1b84: x = 16'h2994; 14'h1b85: x = 16'h2993; 14'h1b86: x = 16'h2992; 14'h1b87: x = 16'h2991; 14'h1b88: x = 16'h2990; 14'h1b89: x = 16'h298f; 14'h1b8a: x = 16'h298e; 14'h1b8b: x = 16'h298d; 14'h1b8c: x = 16'h298c; 14'h1b8d: x = 16'h298c; 14'h1b8e: x = 16'h298b; 14'h1b8f: x = 16'h298a; 14'h1b90: x = 16'h2989; 14'h1b91: x = 16'h2988; 14'h1b92: x = 16'h2987; 14'h1b93: x = 16'h2986; 14'h1b94: x = 16'h2985; 14'h1b95: x = 16'h2984; 14'h1b96: x = 16'h2984; 14'h1b97: x = 16'h2983; 14'h1b98: x = 16'h2982; 14'h1b99: x = 16'h2981; 14'h1b9a: x = 16'h2980; 14'h1b9b: x = 16'h297f; 14'h1b9c: x = 16'h297e; 14'h1b9d: x = 16'h297d; 14'h1b9e: x = 16'h297c; 14'h1b9f: x = 16'h297b; 14'h1ba0: x = 16'h297b; 14'h1ba1: x = 16'h297a; 14'h1ba2: x = 16'h2979; 14'h1ba3: x = 16'h2978; 14'h1ba4: x = 16'h2977; 14'h1ba5: x = 16'h2976; 14'h1ba6: x = 16'h2975; 14'h1ba7: x = 16'h2974; 14'h1ba8: x = 16'h2973; 14'h1ba9: x = 16'h2973; 14'h1baa: x = 16'h2972; 14'h1bab: x = 16'h2971; 14'h1bac: x = 16'h2970; 14'h1bad: x = 16'h296f; 14'h1bae: x = 16'h296e; 14'h1baf: x = 16'h296d; 14'h1bb0: x = 16'h296c; 14'h1bb1: x = 16'h296b; 14'h1bb2: x = 16'h296a; 14'h1bb3: x = 16'h296a; 14'h1bb4: x = 16'h2969; 14'h1bb5: x = 16'h2968; 14'h1bb6: x = 16'h2967; 14'h1bb7: x = 16'h2966; 14'h1bb8: x = 16'h2965; 14'h1bb9: x = 16'h2964; 14'h1bba: x = 16'h2963; 14'h1bbb: x = 16'h2962; 14'h1bbc: x = 16'h2962; 14'h1bbd: x = 16'h2961; 14'h1bbe: x = 16'h2960; 14'h1bbf: x = 16'h295f; 14'h1bc0: x = 16'h295e; 14'h1bc1: x = 16'h295d; 14'h1bc2: x = 16'h295c; 14'h1bc3: x = 16'h295b; 14'h1bc4: x = 16'h295a; 14'h1bc5: x = 16'h295a; 14'h1bc6: x = 16'h2959; 14'h1bc7: x = 16'h2958; 14'h1bc8: x = 16'h2957; 14'h1bc9: x = 16'h2956; 14'h1bca: x = 16'h2955; 14'h1bcb: x = 16'h2954; 14'h1bcc: x = 16'h2953; 14'h1bcd: x = 16'h2952; 14'h1bce: x = 16'h2952; 14'h1bcf: x = 16'h2951; 14'h1bd0: x = 16'h2950; 14'h1bd1: x = 16'h294f; 14'h1bd2: x = 16'h294e; 14'h1bd3: x = 16'h294d; 14'h1bd4: x = 16'h294c; 14'h1bd5: x = 16'h294b; 14'h1bd6: x = 16'h294a; 14'h1bd7: x = 16'h2949; 14'h1bd8: x = 16'h2949; 14'h1bd9: x = 16'h2948; 14'h1bda: x = 16'h2947; 14'h1bdb: x = 16'h2946; 14'h1bdc: x = 16'h2945; 14'h1bdd: x = 16'h2944; 14'h1bde: x = 16'h2943; 14'h1bdf: x = 16'h2942; 14'h1be0: x = 16'h2941; 14'h1be1: x = 16'h2941; 14'h1be2: x = 16'h2940; 14'h1be3: x = 16'h293f; 14'h1be4: x = 16'h293e; 14'h1be5: x = 16'h293d; 14'h1be6: x = 16'h293c; 14'h1be7: x = 16'h293b; 14'h1be8: x = 16'h293a; 14'h1be9: x = 16'h2939; 14'h1bea: x = 16'h2939; 14'h1beb: x = 16'h2938; 14'h1bec: x = 16'h2937; 14'h1bed: x = 16'h2936; 14'h1bee: x = 16'h2935; 14'h1bef: x = 16'h2934; 14'h1bf0: x = 16'h2933; 14'h1bf1: x = 16'h2932; 14'h1bf2: x = 16'h2931; 14'h1bf3: x = 16'h2931; 14'h1bf4: x = 16'h2930; 14'h1bf5: x = 16'h292f; 14'h1bf6: x = 16'h292e; 14'h1bf7: x = 16'h292d; 14'h1bf8: x = 16'h292c; 14'h1bf9: x = 16'h292b; 14'h1bfa: x = 16'h292a; 14'h1bfb: x = 16'h2929; 14'h1bfc: x = 16'h2929; 14'h1bfd: x = 16'h2928; 14'h1bfe: x = 16'h2927; 14'h1bff: x = 16'h2926; 14'h1c00: x = 16'h2925; 14'h1c01: x = 16'h2924; 14'h1c02: x = 16'h2923; 14'h1c03: x = 16'h2922; 14'h1c04: x = 16'h2921; 14'h1c05: x = 16'h2921; 14'h1c06: x = 16'h2920; 14'h1c07: x = 16'h291f; 14'h1c08: x = 16'h291e; 14'h1c09: x = 16'h291d; 14'h1c0a: x = 16'h291c; 14'h1c0b: x = 16'h291b; 14'h1c0c: x = 16'h291a; 14'h1c0d: x = 16'h2919; 14'h1c0e: x = 16'h2919; 14'h1c0f: x = 16'h2918; 14'h1c10: x = 16'h2917; 14'h1c11: x = 16'h2916; 14'h1c12: x = 16'h2915; 14'h1c13: x = 16'h2914; 14'h1c14: x = 16'h2913; 14'h1c15: x = 16'h2912; 14'h1c16: x = 16'h2911; 14'h1c17: x = 16'h2911; 14'h1c18: x = 16'h2910; 14'h1c19: x = 16'h290f; 14'h1c1a: x = 16'h290e; 14'h1c1b: x = 16'h290d; 14'h1c1c: x = 16'h290c; 14'h1c1d: x = 16'h290b; 14'h1c1e: x = 16'h290a; 14'h1c1f: x = 16'h2909; 14'h1c20: x = 16'h2909; 14'h1c21: x = 16'h2908; 14'h1c22: x = 16'h2907; 14'h1c23: x = 16'h2906; 14'h1c24: x = 16'h2905; 14'h1c25: x = 16'h2904; 14'h1c26: x = 16'h2903; 14'h1c27: x = 16'h2902; 14'h1c28: x = 16'h2902; 14'h1c29: x = 16'h2901; 14'h1c2a: x = 16'h2900; 14'h1c2b: x = 16'h28ff; 14'h1c2c: x = 16'h28fe; 14'h1c2d: x = 16'h28fd; 14'h1c2e: x = 16'h28fc; 14'h1c2f: x = 16'h28fb; 14'h1c30: x = 16'h28fa; 14'h1c31: x = 16'h28fa; 14'h1c32: x = 16'h28f9; 14'h1c33: x = 16'h28f8; 14'h1c34: x = 16'h28f7; 14'h1c35: x = 16'h28f6; 14'h1c36: x = 16'h28f5; 14'h1c37: x = 16'h28f4; 14'h1c38: x = 16'h28f3; 14'h1c39: x = 16'h28f2; 14'h1c3a: x = 16'h28f2; 14'h1c3b: x = 16'h28f1; 14'h1c3c: x = 16'h28f0; 14'h1c3d: x = 16'h28ef; 14'h1c3e: x = 16'h28ee; 14'h1c3f: x = 16'h28ed; 14'h1c40: x = 16'h28ec; 14'h1c41: x = 16'h28eb; 14'h1c42: x = 16'h28ea; 14'h1c43: x = 16'h28ea; 14'h1c44: x = 16'h28e9; 14'h1c45: x = 16'h28e8; 14'h1c46: x = 16'h28e7; 14'h1c47: x = 16'h28e6; 14'h1c48: x = 16'h28e5; 14'h1c49: x = 16'h28e4; 14'h1c4a: x = 16'h28e3; 14'h1c4b: x = 16'h28e2; 14'h1c4c: x = 16'h28e2; 14'h1c4d: x = 16'h28e1; 14'h1c4e: x = 16'h28e0; 14'h1c4f: x = 16'h28df; 14'h1c50: x = 16'h28de; 14'h1c51: x = 16'h28dd; 14'h1c52: x = 16'h28dc; 14'h1c53: x = 16'h28db; 14'h1c54: x = 16'h28db; 14'h1c55: x = 16'h28da; 14'h1c56: x = 16'h28d9; 14'h1c57: x = 16'h28d8; 14'h1c58: x = 16'h28d7; 14'h1c59: x = 16'h28d6; 14'h1c5a: x = 16'h28d5; 14'h1c5b: x = 16'h28d4; 14'h1c5c: x = 16'h28d3; 14'h1c5d: x = 16'h28d3; 14'h1c5e: x = 16'h28d2; 14'h1c5f: x = 16'h28d1; 14'h1c60: x = 16'h28d0; 14'h1c61: x = 16'h28cf; 14'h1c62: x = 16'h28ce; 14'h1c63: x = 16'h28cd; 14'h1c64: x = 16'h28cc; 14'h1c65: x = 16'h28cb; 14'h1c66: x = 16'h28cb; 14'h1c67: x = 16'h28ca; 14'h1c68: x = 16'h28c9; 14'h1c69: x = 16'h28c8; 14'h1c6a: x = 16'h28c7; 14'h1c6b: x = 16'h28c6; 14'h1c6c: x = 16'h28c5; 14'h1c6d: x = 16'h28c4; 14'h1c6e: x = 16'h28c4; 14'h1c6f: x = 16'h28c3; 14'h1c70: x = 16'h28c2; 14'h1c71: x = 16'h28c1; 14'h1c72: x = 16'h28c0; 14'h1c73: x = 16'h28bf; 14'h1c74: x = 16'h28be; 14'h1c75: x = 16'h28bd; 14'h1c76: x = 16'h28bc; 14'h1c77: x = 16'h28bc; 14'h1c78: x = 16'h28bb; 14'h1c79: x = 16'h28ba; 14'h1c7a: x = 16'h28b9; 14'h1c7b: x = 16'h28b8; 14'h1c7c: x = 16'h28b7; 14'h1c7d: x = 16'h28b6; 14'h1c7e: x = 16'h28b5; 14'h1c7f: x = 16'h28b5; 14'h1c80: x = 16'h28b4; 14'h1c81: x = 16'h28b3; 14'h1c82: x = 16'h28b2; 14'h1c83: x = 16'h28b1; 14'h1c84: x = 16'h28b0; 14'h1c85: x = 16'h28af; 14'h1c86: x = 16'h28ae; 14'h1c87: x = 16'h28ad; 14'h1c88: x = 16'h28ad; 14'h1c89: x = 16'h28ac; 14'h1c8a: x = 16'h28ab; 14'h1c8b: x = 16'h28aa; 14'h1c8c: x = 16'h28a9; 14'h1c8d: x = 16'h28a8; 14'h1c8e: x = 16'h28a7; 14'h1c8f: x = 16'h28a6; 14'h1c90: x = 16'h28a6; 14'h1c91: x = 16'h28a5; 14'h1c92: x = 16'h28a4; 14'h1c93: x = 16'h28a3; 14'h1c94: x = 16'h28a2; 14'h1c95: x = 16'h28a1; 14'h1c96: x = 16'h28a0; 14'h1c97: x = 16'h289f; 14'h1c98: x = 16'h289e; 14'h1c99: x = 16'h289e; 14'h1c9a: x = 16'h289d; 14'h1c9b: x = 16'h289c; 14'h1c9c: x = 16'h289b; 14'h1c9d: x = 16'h289a; 14'h1c9e: x = 16'h2899; 14'h1c9f: x = 16'h2898; 14'h1ca0: x = 16'h2897; 14'h1ca1: x = 16'h2897; 14'h1ca2: x = 16'h2896; 14'h1ca3: x = 16'h2895; 14'h1ca4: x = 16'h2894; 14'h1ca5: x = 16'h2893; 14'h1ca6: x = 16'h2892; 14'h1ca7: x = 16'h2891; 14'h1ca8: x = 16'h2890; 14'h1ca9: x = 16'h288f; 14'h1caa: x = 16'h288f; 14'h1cab: x = 16'h288e; 14'h1cac: x = 16'h288d; 14'h1cad: x = 16'h288c; 14'h1cae: x = 16'h288b; 14'h1caf: x = 16'h288a; 14'h1cb0: x = 16'h2889; 14'h1cb1: x = 16'h2888; 14'h1cb2: x = 16'h2888; 14'h1cb3: x = 16'h2887; 14'h1cb4: x = 16'h2886; 14'h1cb5: x = 16'h2885; 14'h1cb6: x = 16'h2884; 14'h1cb7: x = 16'h2883; 14'h1cb8: x = 16'h2882; 14'h1cb9: x = 16'h2881; 14'h1cba: x = 16'h2881; 14'h1cbb: x = 16'h2880; 14'h1cbc: x = 16'h287f; 14'h1cbd: x = 16'h287e; 14'h1cbe: x = 16'h287d; 14'h1cbf: x = 16'h287c; 14'h1cc0: x = 16'h287b; 14'h1cc1: x = 16'h287a; 14'h1cc2: x = 16'h2879; 14'h1cc3: x = 16'h2879; 14'h1cc4: x = 16'h2878; 14'h1cc5: x = 16'h2877; 14'h1cc6: x = 16'h2876; 14'h1cc7: x = 16'h2875; 14'h1cc8: x = 16'h2874; 14'h1cc9: x = 16'h2873; 14'h1cca: x = 16'h2872; 14'h1ccb: x = 16'h2872; 14'h1ccc: x = 16'h2871; 14'h1ccd: x = 16'h2870; 14'h1cce: x = 16'h286f; 14'h1ccf: x = 16'h286e; 14'h1cd0: x = 16'h286d; 14'h1cd1: x = 16'h286c; 14'h1cd2: x = 16'h286b; 14'h1cd3: x = 16'h286b; 14'h1cd4: x = 16'h286a; 14'h1cd5: x = 16'h2869; 14'h1cd6: x = 16'h2868; 14'h1cd7: x = 16'h2867; 14'h1cd8: x = 16'h2866; 14'h1cd9: x = 16'h2865; 14'h1cda: x = 16'h2864; 14'h1cdb: x = 16'h2864; 14'h1cdc: x = 16'h2863; 14'h1cdd: x = 16'h2862; 14'h1cde: x = 16'h2861; 14'h1cdf: x = 16'h2860; 14'h1ce0: x = 16'h285f; 14'h1ce1: x = 16'h285e; 14'h1ce2: x = 16'h285d; 14'h1ce3: x = 16'h285c; 14'h1ce4: x = 16'h285c; 14'h1ce5: x = 16'h285b; 14'h1ce6: x = 16'h285a; 14'h1ce7: x = 16'h2859; 14'h1ce8: x = 16'h2858; 14'h1ce9: x = 16'h2857; 14'h1cea: x = 16'h2856; 14'h1ceb: x = 16'h2855; 14'h1cec: x = 16'h2855; 14'h1ced: x = 16'h2854; 14'h1cee: x = 16'h2853; 14'h1cef: x = 16'h2852; 14'h1cf0: x = 16'h2851; 14'h1cf1: x = 16'h2850; 14'h1cf2: x = 16'h284f; 14'h1cf3: x = 16'h284e; 14'h1cf4: x = 16'h284e; 14'h1cf5: x = 16'h284d; 14'h1cf6: x = 16'h284c; 14'h1cf7: x = 16'h284b; 14'h1cf8: x = 16'h284a; 14'h1cf9: x = 16'h2849; 14'h1cfa: x = 16'h2848; 14'h1cfb: x = 16'h2847; 14'h1cfc: x = 16'h2847; 14'h1cfd: x = 16'h2846; 14'h1cfe: x = 16'h2845; 14'h1cff: x = 16'h2844; 14'h1d00: x = 16'h2843; 14'h1d01: x = 16'h2842; 14'h1d02: x = 16'h2841; 14'h1d03: x = 16'h2840; 14'h1d04: x = 16'h2840; 14'h1d05: x = 16'h283f; 14'h1d06: x = 16'h283e; 14'h1d07: x = 16'h283d; 14'h1d08: x = 16'h283c; 14'h1d09: x = 16'h283b; 14'h1d0a: x = 16'h283a; 14'h1d0b: x = 16'h2839; 14'h1d0c: x = 16'h2839; 14'h1d0d: x = 16'h2838; 14'h1d0e: x = 16'h2837; 14'h1d0f: x = 16'h2836; 14'h1d10: x = 16'h2835; 14'h1d11: x = 16'h2834; 14'h1d12: x = 16'h2833; 14'h1d13: x = 16'h2832; 14'h1d14: x = 16'h2831; 14'h1d15: x = 16'h2831; 14'h1d16: x = 16'h2830; 14'h1d17: x = 16'h282f; 14'h1d18: x = 16'h282e; 14'h1d19: x = 16'h282d; 14'h1d1a: x = 16'h282c; 14'h1d1b: x = 16'h282b; 14'h1d1c: x = 16'h282a; 14'h1d1d: x = 16'h282a; 14'h1d1e: x = 16'h2829; 14'h1d1f: x = 16'h2828; 14'h1d20: x = 16'h2827; 14'h1d21: x = 16'h2826; 14'h1d22: x = 16'h2825; 14'h1d23: x = 16'h2824; 14'h1d24: x = 16'h2823; 14'h1d25: x = 16'h2823; 14'h1d26: x = 16'h2822; 14'h1d27: x = 16'h2821; 14'h1d28: x = 16'h2820; 14'h1d29: x = 16'h281f; 14'h1d2a: x = 16'h281e; 14'h1d2b: x = 16'h281d; 14'h1d2c: x = 16'h281c; 14'h1d2d: x = 16'h281c; 14'h1d2e: x = 16'h281b; 14'h1d2f: x = 16'h281a; 14'h1d30: x = 16'h2819; 14'h1d31: x = 16'h2818; 14'h1d32: x = 16'h2817; 14'h1d33: x = 16'h2816; 14'h1d34: x = 16'h2815; 14'h1d35: x = 16'h2815; 14'h1d36: x = 16'h2814; 14'h1d37: x = 16'h2813; 14'h1d38: x = 16'h2812; 14'h1d39: x = 16'h2811; 14'h1d3a: x = 16'h2810; 14'h1d3b: x = 16'h280f; 14'h1d3c: x = 16'h280e; 14'h1d3d: x = 16'h280e; 14'h1d3e: x = 16'h280d; 14'h1d3f: x = 16'h280c; 14'h1d40: x = 16'h280b; 14'h1d41: x = 16'h280a; 14'h1d42: x = 16'h2809; 14'h1d43: x = 16'h2808; 14'h1d44: x = 16'h2807; 14'h1d45: x = 16'h2807; 14'h1d46: x = 16'h2806; 14'h1d47: x = 16'h2805; 14'h1d48: x = 16'h2804; 14'h1d49: x = 16'h2803; 14'h1d4a: x = 16'h2802; 14'h1d4b: x = 16'h2801; 14'h1d4c: x = 16'h2800; 14'h1d4d: x = 16'h2800; 14'h1d4e: x = 16'h27ff; 14'h1d4f: x = 16'h27fe; 14'h1d50: x = 16'h27fd; 14'h1d51: x = 16'h27fc; 14'h1d52: x = 16'h27fb; 14'h1d53: x = 16'h27fa; 14'h1d54: x = 16'h27fa; 14'h1d55: x = 16'h27f9; 14'h1d56: x = 16'h27f8; 14'h1d57: x = 16'h27f7; 14'h1d58: x = 16'h27f6; 14'h1d59: x = 16'h27f5; 14'h1d5a: x = 16'h27f4; 14'h1d5b: x = 16'h27f3; 14'h1d5c: x = 16'h27f3; 14'h1d5d: x = 16'h27f2; 14'h1d5e: x = 16'h27f1; 14'h1d5f: x = 16'h27f0; 14'h1d60: x = 16'h27ef; 14'h1d61: x = 16'h27ee; 14'h1d62: x = 16'h27ed; 14'h1d63: x = 16'h27ec; 14'h1d64: x = 16'h27ec; 14'h1d65: x = 16'h27eb; 14'h1d66: x = 16'h27ea; 14'h1d67: x = 16'h27e9; 14'h1d68: x = 16'h27e8; 14'h1d69: x = 16'h27e7; 14'h1d6a: x = 16'h27e6; 14'h1d6b: x = 16'h27e5; 14'h1d6c: x = 16'h27e5; 14'h1d6d: x = 16'h27e4; 14'h1d6e: x = 16'h27e3; 14'h1d6f: x = 16'h27e2; 14'h1d70: x = 16'h27e1; 14'h1d71: x = 16'h27e0; 14'h1d72: x = 16'h27df; 14'h1d73: x = 16'h27de; 14'h1d74: x = 16'h27de; 14'h1d75: x = 16'h27dd; 14'h1d76: x = 16'h27dc; 14'h1d77: x = 16'h27db; 14'h1d78: x = 16'h27da; 14'h1d79: x = 16'h27d9; 14'h1d7a: x = 16'h27d8; 14'h1d7b: x = 16'h27d7; 14'h1d7c: x = 16'h27d7; 14'h1d7d: x = 16'h27d6; 14'h1d7e: x = 16'h27d5; 14'h1d7f: x = 16'h27d4; 14'h1d80: x = 16'h27d3; 14'h1d81: x = 16'h27d2; 14'h1d82: x = 16'h27d1; 14'h1d83: x = 16'h27d1; 14'h1d84: x = 16'h27d0; 14'h1d85: x = 16'h27cf; 14'h1d86: x = 16'h27ce; 14'h1d87: x = 16'h27cd; 14'h1d88: x = 16'h27cc; 14'h1d89: x = 16'h27cb; 14'h1d8a: x = 16'h27ca; 14'h1d8b: x = 16'h27ca; 14'h1d8c: x = 16'h27c9; 14'h1d8d: x = 16'h27c8; 14'h1d8e: x = 16'h27c7; 14'h1d8f: x = 16'h27c6; 14'h1d90: x = 16'h27c5; 14'h1d91: x = 16'h27c4; 14'h1d92: x = 16'h27c3; 14'h1d93: x = 16'h27c3; 14'h1d94: x = 16'h27c2; 14'h1d95: x = 16'h27c1; 14'h1d96: x = 16'h27c0; 14'h1d97: x = 16'h27bf; 14'h1d98: x = 16'h27be; 14'h1d99: x = 16'h27bd; 14'h1d9a: x = 16'h27bc; 14'h1d9b: x = 16'h27bc; 14'h1d9c: x = 16'h27bb; 14'h1d9d: x = 16'h27ba; 14'h1d9e: x = 16'h27b9; 14'h1d9f: x = 16'h27b8; 14'h1da0: x = 16'h27b7; 14'h1da1: x = 16'h27b6; 14'h1da2: x = 16'h27b6; 14'h1da3: x = 16'h27b5; 14'h1da4: x = 16'h27b4; 14'h1da5: x = 16'h27b3; 14'h1da6: x = 16'h27b2; 14'h1da7: x = 16'h27b1; 14'h1da8: x = 16'h27b0; 14'h1da9: x = 16'h27af; 14'h1daa: x = 16'h27af; 14'h1dab: x = 16'h27ae; 14'h1dac: x = 16'h27ad; 14'h1dad: x = 16'h27ac; 14'h1dae: x = 16'h27ab; 14'h1daf: x = 16'h27aa; 14'h1db0: x = 16'h27a9; 14'h1db1: x = 16'h27a8; 14'h1db2: x = 16'h27a8; 14'h1db3: x = 16'h27a7; 14'h1db4: x = 16'h27a6; 14'h1db5: x = 16'h27a5; 14'h1db6: x = 16'h27a4; 14'h1db7: x = 16'h27a3; 14'h1db8: x = 16'h27a2; 14'h1db9: x = 16'h27a2; 14'h1dba: x = 16'h27a1; 14'h1dbb: x = 16'h27a0; 14'h1dbc: x = 16'h279f; 14'h1dbd: x = 16'h279e; 14'h1dbe: x = 16'h279d; 14'h1dbf: x = 16'h279c; 14'h1dc0: x = 16'h279b; 14'h1dc1: x = 16'h279b; 14'h1dc2: x = 16'h279a; 14'h1dc3: x = 16'h2799; 14'h1dc4: x = 16'h2798; 14'h1dc5: x = 16'h2797; 14'h1dc6: x = 16'h2796; 14'h1dc7: x = 16'h2795; 14'h1dc8: x = 16'h2794; 14'h1dc9: x = 16'h2794; 14'h1dca: x = 16'h2793; 14'h1dcb: x = 16'h2792; 14'h1dcc: x = 16'h2791; 14'h1dcd: x = 16'h2790; 14'h1dce: x = 16'h278f; 14'h1dcf: x = 16'h278e; 14'h1dd0: x = 16'h278e; 14'h1dd1: x = 16'h278d; 14'h1dd2: x = 16'h278c; 14'h1dd3: x = 16'h278b; 14'h1dd4: x = 16'h278a; 14'h1dd5: x = 16'h2789; 14'h1dd6: x = 16'h2788; 14'h1dd7: x = 16'h2787; 14'h1dd8: x = 16'h2787; 14'h1dd9: x = 16'h2786; 14'h1dda: x = 16'h2785; 14'h1ddb: x = 16'h2784; 14'h1ddc: x = 16'h2783; 14'h1ddd: x = 16'h2782; 14'h1dde: x = 16'h2781; 14'h1ddf: x = 16'h2781; 14'h1de0: x = 16'h2780; 14'h1de1: x = 16'h277f; 14'h1de2: x = 16'h277e; 14'h1de3: x = 16'h277d; 14'h1de4: x = 16'h277c; 14'h1de5: x = 16'h277b; 14'h1de6: x = 16'h277a; 14'h1de7: x = 16'h277a; 14'h1de8: x = 16'h2779; 14'h1de9: x = 16'h2778; 14'h1dea: x = 16'h2777; 14'h1deb: x = 16'h2776; 14'h1dec: x = 16'h2775; 14'h1ded: x = 16'h2774; 14'h1dee: x = 16'h2773; 14'h1def: x = 16'h2773; 14'h1df0: x = 16'h2772; 14'h1df1: x = 16'h2771; 14'h1df2: x = 16'h2770; 14'h1df3: x = 16'h276f; 14'h1df4: x = 16'h276e; 14'h1df5: x = 16'h276d; 14'h1df6: x = 16'h276d; 14'h1df7: x = 16'h276c; 14'h1df8: x = 16'h276b; 14'h1df9: x = 16'h276a; 14'h1dfa: x = 16'h2769; 14'h1dfb: x = 16'h2768; 14'h1dfc: x = 16'h2767; 14'h1dfd: x = 16'h2766; 14'h1dfe: x = 16'h2766; 14'h1dff: x = 16'h2765; 14'h1e00: x = 16'h2764; 14'h1e01: x = 16'h2763; 14'h1e02: x = 16'h2762; 14'h1e03: x = 16'h2761; 14'h1e04: x = 16'h2760; 14'h1e05: x = 16'h2760; 14'h1e06: x = 16'h275f; 14'h1e07: x = 16'h275e; 14'h1e08: x = 16'h275d; 14'h1e09: x = 16'h275c; 14'h1e0a: x = 16'h275b; 14'h1e0b: x = 16'h275a; 14'h1e0c: x = 16'h2759; 14'h1e0d: x = 16'h2759; 14'h1e0e: x = 16'h2758; 14'h1e0f: x = 16'h2757; 14'h1e10: x = 16'h2756; 14'h1e11: x = 16'h2755; 14'h1e12: x = 16'h2754; 14'h1e13: x = 16'h2753; 14'h1e14: x = 16'h2753; 14'h1e15: x = 16'h2752; 14'h1e16: x = 16'h2751; 14'h1e17: x = 16'h2750; 14'h1e18: x = 16'h274f; 14'h1e19: x = 16'h274e; 14'h1e1a: x = 16'h274d; 14'h1e1b: x = 16'h274d; 14'h1e1c: x = 16'h274c; 14'h1e1d: x = 16'h274b; 14'h1e1e: x = 16'h274a; 14'h1e1f: x = 16'h2749; 14'h1e20: x = 16'h2748; 14'h1e21: x = 16'h2747; 14'h1e22: x = 16'h2746; 14'h1e23: x = 16'h2746; 14'h1e24: x = 16'h2745; 14'h1e25: x = 16'h2744; 14'h1e26: x = 16'h2743; 14'h1e27: x = 16'h2742; 14'h1e28: x = 16'h2741; 14'h1e29: x = 16'h2740; 14'h1e2a: x = 16'h2740; 14'h1e2b: x = 16'h273f; 14'h1e2c: x = 16'h273e; 14'h1e2d: x = 16'h273d; 14'h1e2e: x = 16'h273c; 14'h1e2f: x = 16'h273b; 14'h1e30: x = 16'h273a; 14'h1e31: x = 16'h2739; 14'h1e32: x = 16'h2739; 14'h1e33: x = 16'h2738; 14'h1e34: x = 16'h2737; 14'h1e35: x = 16'h2736; 14'h1e36: x = 16'h2735; 14'h1e37: x = 16'h2734; 14'h1e38: x = 16'h2733; 14'h1e39: x = 16'h2733; 14'h1e3a: x = 16'h2732; 14'h1e3b: x = 16'h2731; 14'h1e3c: x = 16'h2730; 14'h1e3d: x = 16'h272f; 14'h1e3e: x = 16'h272e; 14'h1e3f: x = 16'h272d; 14'h1e40: x = 16'h272d; 14'h1e41: x = 16'h272c; 14'h1e42: x = 16'h272b; 14'h1e43: x = 16'h272a; 14'h1e44: x = 16'h2729; 14'h1e45: x = 16'h2728; 14'h1e46: x = 16'h2727; 14'h1e47: x = 16'h2726; 14'h1e48: x = 16'h2726; 14'h1e49: x = 16'h2725; 14'h1e4a: x = 16'h2724; 14'h1e4b: x = 16'h2723; 14'h1e4c: x = 16'h2722; 14'h1e4d: x = 16'h2721; 14'h1e4e: x = 16'h2720; 14'h1e4f: x = 16'h2720; 14'h1e50: x = 16'h271f; 14'h1e51: x = 16'h271e; 14'h1e52: x = 16'h271d; 14'h1e53: x = 16'h271c; 14'h1e54: x = 16'h271b; 14'h1e55: x = 16'h271a; 14'h1e56: x = 16'h271a; 14'h1e57: x = 16'h2719; 14'h1e58: x = 16'h2718; 14'h1e59: x = 16'h2717; 14'h1e5a: x = 16'h2716; 14'h1e5b: x = 16'h2715; 14'h1e5c: x = 16'h2714; 14'h1e5d: x = 16'h2713; 14'h1e5e: x = 16'h2713; 14'h1e5f: x = 16'h2712; 14'h1e60: x = 16'h2711; 14'h1e61: x = 16'h2710; 14'h1e62: x = 16'h270f; 14'h1e63: x = 16'h270e; 14'h1e64: x = 16'h270d; 14'h1e65: x = 16'h270d; 14'h1e66: x = 16'h270c; 14'h1e67: x = 16'h270b; 14'h1e68: x = 16'h270a; 14'h1e69: x = 16'h2709; 14'h1e6a: x = 16'h2708; 14'h1e6b: x = 16'h2707; 14'h1e6c: x = 16'h2707; 14'h1e6d: x = 16'h2706; 14'h1e6e: x = 16'h2705; 14'h1e6f: x = 16'h2704; 14'h1e70: x = 16'h2703; 14'h1e71: x = 16'h2702; 14'h1e72: x = 16'h2701; 14'h1e73: x = 16'h2700; 14'h1e74: x = 16'h2700; 14'h1e75: x = 16'h26ff; 14'h1e76: x = 16'h26fe; 14'h1e77: x = 16'h26fd; 14'h1e78: x = 16'h26fc; 14'h1e79: x = 16'h26fb; 14'h1e7a: x = 16'h26fa; 14'h1e7b: x = 16'h26fa; 14'h1e7c: x = 16'h26f9; 14'h1e7d: x = 16'h26f8; 14'h1e7e: x = 16'h26f7; 14'h1e7f: x = 16'h26f6; 14'h1e80: x = 16'h26f5; 14'h1e81: x = 16'h26f4; 14'h1e82: x = 16'h26f4; 14'h1e83: x = 16'h26f3; 14'h1e84: x = 16'h26f2; 14'h1e85: x = 16'h26f1; 14'h1e86: x = 16'h26f0; 14'h1e87: x = 16'h26ef; 14'h1e88: x = 16'h26ee; 14'h1e89: x = 16'h26ee; 14'h1e8a: x = 16'h26ed; 14'h1e8b: x = 16'h26ec; 14'h1e8c: x = 16'h26eb; 14'h1e8d: x = 16'h26ea; 14'h1e8e: x = 16'h26e9; 14'h1e8f: x = 16'h26e8; 14'h1e90: x = 16'h26e7; 14'h1e91: x = 16'h26e7; 14'h1e92: x = 16'h26e6; 14'h1e93: x = 16'h26e5; 14'h1e94: x = 16'h26e4; 14'h1e95: x = 16'h26e3; 14'h1e96: x = 16'h26e2; 14'h1e97: x = 16'h26e1; 14'h1e98: x = 16'h26e1; 14'h1e99: x = 16'h26e0; 14'h1e9a: x = 16'h26df; 14'h1e9b: x = 16'h26de; 14'h1e9c: x = 16'h26dd; 14'h1e9d: x = 16'h26dc; 14'h1e9e: x = 16'h26db; 14'h1e9f: x = 16'h26db; 14'h1ea0: x = 16'h26da; 14'h1ea1: x = 16'h26d9; 14'h1ea2: x = 16'h26d8; 14'h1ea3: x = 16'h26d7; 14'h1ea4: x = 16'h26d6; 14'h1ea5: x = 16'h26d5; 14'h1ea6: x = 16'h26d5; 14'h1ea7: x = 16'h26d4; 14'h1ea8: x = 16'h26d3; 14'h1ea9: x = 16'h26d2; 14'h1eaa: x = 16'h26d1; 14'h1eab: x = 16'h26d0; 14'h1eac: x = 16'h26cf; 14'h1ead: x = 16'h26cf; 14'h1eae: x = 16'h26ce; 14'h1eaf: x = 16'h26cd; 14'h1eb0: x = 16'h26cc; 14'h1eb1: x = 16'h26cb; 14'h1eb2: x = 16'h26ca; 14'h1eb3: x = 16'h26c9; 14'h1eb4: x = 16'h26c9; 14'h1eb5: x = 16'h26c8; 14'h1eb6: x = 16'h26c7; 14'h1eb7: x = 16'h26c6; 14'h1eb8: x = 16'h26c5; 14'h1eb9: x = 16'h26c4; 14'h1eba: x = 16'h26c3; 14'h1ebb: x = 16'h26c3; 14'h1ebc: x = 16'h26c2; 14'h1ebd: x = 16'h26c1; 14'h1ebe: x = 16'h26c0; 14'h1ebf: x = 16'h26bf; 14'h1ec0: x = 16'h26be; 14'h1ec1: x = 16'h26bd; 14'h1ec2: x = 16'h26bc; 14'h1ec3: x = 16'h26bc; 14'h1ec4: x = 16'h26bb; 14'h1ec5: x = 16'h26ba; 14'h1ec6: x = 16'h26b9; 14'h1ec7: x = 16'h26b8; 14'h1ec8: x = 16'h26b7; 14'h1ec9: x = 16'h26b6; 14'h1eca: x = 16'h26b6; 14'h1ecb: x = 16'h26b5; 14'h1ecc: x = 16'h26b4; 14'h1ecd: x = 16'h26b3; 14'h1ece: x = 16'h26b2; 14'h1ecf: x = 16'h26b1; 14'h1ed0: x = 16'h26b0; 14'h1ed1: x = 16'h26b0; 14'h1ed2: x = 16'h26af; 14'h1ed3: x = 16'h26ae; 14'h1ed4: x = 16'h26ad; 14'h1ed5: x = 16'h26ac; 14'h1ed6: x = 16'h26ab; 14'h1ed7: x = 16'h26aa; 14'h1ed8: x = 16'h26aa; 14'h1ed9: x = 16'h26a9; 14'h1eda: x = 16'h26a8; 14'h1edb: x = 16'h26a7; 14'h1edc: x = 16'h26a6; 14'h1edd: x = 16'h26a5; 14'h1ede: x = 16'h26a4; 14'h1edf: x = 16'h26a4; 14'h1ee0: x = 16'h26a3; 14'h1ee1: x = 16'h26a2; 14'h1ee2: x = 16'h26a1; 14'h1ee3: x = 16'h26a0; 14'h1ee4: x = 16'h269f; 14'h1ee5: x = 16'h269e; 14'h1ee6: x = 16'h269e; 14'h1ee7: x = 16'h269d; 14'h1ee8: x = 16'h269c; 14'h1ee9: x = 16'h269b; 14'h1eea: x = 16'h269a; 14'h1eeb: x = 16'h2699; 14'h1eec: x = 16'h2698; 14'h1eed: x = 16'h2698; 14'h1eee: x = 16'h2697; 14'h1eef: x = 16'h2696; 14'h1ef0: x = 16'h2695; 14'h1ef1: x = 16'h2694; 14'h1ef2: x = 16'h2693; 14'h1ef3: x = 16'h2692; 14'h1ef4: x = 16'h2692; 14'h1ef5: x = 16'h2691; 14'h1ef6: x = 16'h2690; 14'h1ef7: x = 16'h268f; 14'h1ef8: x = 16'h268e; 14'h1ef9: x = 16'h268d; 14'h1efa: x = 16'h268c; 14'h1efb: x = 16'h268c; 14'h1efc: x = 16'h268b; 14'h1efd: x = 16'h268a; 14'h1efe: x = 16'h2689; 14'h1eff: x = 16'h2688; 14'h1f00: x = 16'h2687; 14'h1f01: x = 16'h2686; 14'h1f02: x = 16'h2686; 14'h1f03: x = 16'h2685; 14'h1f04: x = 16'h2684; 14'h1f05: x = 16'h2683; 14'h1f06: x = 16'h2682; 14'h1f07: x = 16'h2681; 14'h1f08: x = 16'h2680; 14'h1f09: x = 16'h2680; 14'h1f0a: x = 16'h267f; 14'h1f0b: x = 16'h267e; 14'h1f0c: x = 16'h267d; 14'h1f0d: x = 16'h267c; 14'h1f0e: x = 16'h267b; 14'h1f0f: x = 16'h267a; 14'h1f10: x = 16'h267a; 14'h1f11: x = 16'h2679; 14'h1f12: x = 16'h2678; 14'h1f13: x = 16'h2677; 14'h1f14: x = 16'h2676; 14'h1f15: x = 16'h2675; 14'h1f16: x = 16'h2674; 14'h1f17: x = 16'h2674; 14'h1f18: x = 16'h2673; 14'h1f19: x = 16'h2672; 14'h1f1a: x = 16'h2671; 14'h1f1b: x = 16'h2670; 14'h1f1c: x = 16'h266f; 14'h1f1d: x = 16'h266e; 14'h1f1e: x = 16'h266e; 14'h1f1f: x = 16'h266d; 14'h1f20: x = 16'h266c; 14'h1f21: x = 16'h266b; 14'h1f22: x = 16'h266a; 14'h1f23: x = 16'h2669; 14'h1f24: x = 16'h2668; 14'h1f25: x = 16'h2668; 14'h1f26: x = 16'h2667; 14'h1f27: x = 16'h2666; 14'h1f28: x = 16'h2665; 14'h1f29: x = 16'h2664; 14'h1f2a: x = 16'h2663; 14'h1f2b: x = 16'h2662; 14'h1f2c: x = 16'h2662; 14'h1f2d: x = 16'h2661; 14'h1f2e: x = 16'h2660; 14'h1f2f: x = 16'h265f; 14'h1f30: x = 16'h265e; 14'h1f31: x = 16'h265d; 14'h1f32: x = 16'h265c; 14'h1f33: x = 16'h265c; 14'h1f34: x = 16'h265b; 14'h1f35: x = 16'h265a; 14'h1f36: x = 16'h2659; 14'h1f37: x = 16'h2658; 14'h1f38: x = 16'h2657; 14'h1f39: x = 16'h2656; 14'h1f3a: x = 16'h2656; 14'h1f3b: x = 16'h2655; 14'h1f3c: x = 16'h2654; 14'h1f3d: x = 16'h2653; 14'h1f3e: x = 16'h2652; 14'h1f3f: x = 16'h2651; 14'h1f40: x = 16'h2650; 14'h1f41: x = 16'h2650; 14'h1f42: x = 16'h264f; 14'h1f43: x = 16'h264e; 14'h1f44: x = 16'h264d; 14'h1f45: x = 16'h264c; 14'h1f46: x = 16'h264b; 14'h1f47: x = 16'h264a; 14'h1f48: x = 16'h264a; 14'h1f49: x = 16'h2649; 14'h1f4a: x = 16'h2648; 14'h1f4b: x = 16'h2647; 14'h1f4c: x = 16'h2646; 14'h1f4d: x = 16'h2645; 14'h1f4e: x = 16'h2644; 14'h1f4f: x = 16'h2644; 14'h1f50: x = 16'h2643; 14'h1f51: x = 16'h2642; 14'h1f52: x = 16'h2641; 14'h1f53: x = 16'h2640; 14'h1f54: x = 16'h263f; 14'h1f55: x = 16'h263f; 14'h1f56: x = 16'h263e; 14'h1f57: x = 16'h263d; 14'h1f58: x = 16'h263c; 14'h1f59: x = 16'h263b; 14'h1f5a: x = 16'h263a; 14'h1f5b: x = 16'h2639; 14'h1f5c: x = 16'h2639; 14'h1f5d: x = 16'h2638; 14'h1f5e: x = 16'h2637; 14'h1f5f: x = 16'h2636; 14'h1f60: x = 16'h2635; 14'h1f61: x = 16'h2634; 14'h1f62: x = 16'h2633; 14'h1f63: x = 16'h2633; 14'h1f64: x = 16'h2632; 14'h1f65: x = 16'h2631; 14'h1f66: x = 16'h2630; 14'h1f67: x = 16'h262f; 14'h1f68: x = 16'h262e; 14'h1f69: x = 16'h262d; 14'h1f6a: x = 16'h262d; 14'h1f6b: x = 16'h262c; 14'h1f6c: x = 16'h262b; 14'h1f6d: x = 16'h262a; 14'h1f6e: x = 16'h2629; 14'h1f6f: x = 16'h2628; 14'h1f70: x = 16'h2627; 14'h1f71: x = 16'h2627; 14'h1f72: x = 16'h2626; 14'h1f73: x = 16'h2625; 14'h1f74: x = 16'h2624; 14'h1f75: x = 16'h2623; 14'h1f76: x = 16'h2622; 14'h1f77: x = 16'h2621; 14'h1f78: x = 16'h2621; 14'h1f79: x = 16'h2620; 14'h1f7a: x = 16'h261f; 14'h1f7b: x = 16'h261e; 14'h1f7c: x = 16'h261d; 14'h1f7d: x = 16'h261c; 14'h1f7e: x = 16'h261c; 14'h1f7f: x = 16'h261b; 14'h1f80: x = 16'h261a; 14'h1f81: x = 16'h2619; 14'h1f82: x = 16'h2618; 14'h1f83: x = 16'h2617; 14'h1f84: x = 16'h2616; 14'h1f85: x = 16'h2616; 14'h1f86: x = 16'h2615; 14'h1f87: x = 16'h2614; 14'h1f88: x = 16'h2613; 14'h1f89: x = 16'h2612; 14'h1f8a: x = 16'h2611; 14'h1f8b: x = 16'h2610; 14'h1f8c: x = 16'h2610; 14'h1f8d: x = 16'h260f; 14'h1f8e: x = 16'h260e; 14'h1f8f: x = 16'h260d; 14'h1f90: x = 16'h260c; 14'h1f91: x = 16'h260b; 14'h1f92: x = 16'h260a; 14'h1f93: x = 16'h260a; 14'h1f94: x = 16'h2609; 14'h1f95: x = 16'h2608; 14'h1f96: x = 16'h2607; 14'h1f97: x = 16'h2606; 14'h1f98: x = 16'h2605; 14'h1f99: x = 16'h2604; 14'h1f9a: x = 16'h2604; 14'h1f9b: x = 16'h2603; 14'h1f9c: x = 16'h2602; 14'h1f9d: x = 16'h2601; 14'h1f9e: x = 16'h2600; 14'h1f9f: x = 16'h25ff; 14'h1fa0: x = 16'h25ff; 14'h1fa1: x = 16'h25fe; 14'h1fa2: x = 16'h25fd; 14'h1fa3: x = 16'h25fc; 14'h1fa4: x = 16'h25fb; 14'h1fa5: x = 16'h25fa; 14'h1fa6: x = 16'h25f9; 14'h1fa7: x = 16'h25f9; 14'h1fa8: x = 16'h25f8; 14'h1fa9: x = 16'h25f7; 14'h1faa: x = 16'h25f6; 14'h1fab: x = 16'h25f5; 14'h1fac: x = 16'h25f4; 14'h1fad: x = 16'h25f3; 14'h1fae: x = 16'h25f3; 14'h1faf: x = 16'h25f2; 14'h1fb0: x = 16'h25f1; 14'h1fb1: x = 16'h25f0; 14'h1fb2: x = 16'h25ef; 14'h1fb3: x = 16'h25ee; 14'h1fb4: x = 16'h25ed; 14'h1fb5: x = 16'h25ed; 14'h1fb6: x = 16'h25ec; 14'h1fb7: x = 16'h25eb; 14'h1fb8: x = 16'h25ea; 14'h1fb9: x = 16'h25e9; 14'h1fba: x = 16'h25e8; 14'h1fbb: x = 16'h25e8; 14'h1fbc: x = 16'h25e7; 14'h1fbd: x = 16'h25e6; 14'h1fbe: x = 16'h25e5; 14'h1fbf: x = 16'h25e4; 14'h1fc0: x = 16'h25e3; 14'h1fc1: x = 16'h25e2; 14'h1fc2: x = 16'h25e2; 14'h1fc3: x = 16'h25e1; 14'h1fc4: x = 16'h25e0; 14'h1fc5: x = 16'h25df; 14'h1fc6: x = 16'h25de; 14'h1fc7: x = 16'h25dd; 14'h1fc8: x = 16'h25dc; 14'h1fc9: x = 16'h25dc; 14'h1fca: x = 16'h25db; 14'h1fcb: x = 16'h25da; 14'h1fcc: x = 16'h25d9; 14'h1fcd: x = 16'h25d8; 14'h1fce: x = 16'h25d7; 14'h1fcf: x = 16'h25d6; 14'h1fd0: x = 16'h25d6; 14'h1fd1: x = 16'h25d5; 14'h1fd2: x = 16'h25d4; 14'h1fd3: x = 16'h25d3; 14'h1fd4: x = 16'h25d2; 14'h1fd5: x = 16'h25d1; 14'h1fd6: x = 16'h25d1; 14'h1fd7: x = 16'h25d0; 14'h1fd8: x = 16'h25cf; 14'h1fd9: x = 16'h25ce; 14'h1fda: x = 16'h25cd; 14'h1fdb: x = 16'h25cc; 14'h1fdc: x = 16'h25cb; 14'h1fdd: x = 16'h25cb; 14'h1fde: x = 16'h25ca; 14'h1fdf: x = 16'h25c9; 14'h1fe0: x = 16'h25c8; 14'h1fe1: x = 16'h25c7; 14'h1fe2: x = 16'h25c6; 14'h1fe3: x = 16'h25c5; 14'h1fe4: x = 16'h25c5; 14'h1fe5: x = 16'h25c4; 14'h1fe6: x = 16'h25c3; 14'h1fe7: x = 16'h25c2; 14'h1fe8: x = 16'h25c1; 14'h1fe9: x = 16'h25c0; 14'h1fea: x = 16'h25c0; 14'h1feb: x = 16'h25bf; 14'h1fec: x = 16'h25be; 14'h1fed: x = 16'h25bd; 14'h1fee: x = 16'h25bc; 14'h1fef: x = 16'h25bb; 14'h1ff0: x = 16'h25ba; 14'h1ff1: x = 16'h25ba; 14'h1ff2: x = 16'h25b9; 14'h1ff3: x = 16'h25b8; 14'h1ff4: x = 16'h25b7; 14'h1ff5: x = 16'h25b6; 14'h1ff6: x = 16'h25b5; 14'h1ff7: x = 16'h25b4; 14'h1ff8: x = 16'h25b4; 14'h1ff9: x = 16'h25b3; 14'h1ffa: x = 16'h25b2; 14'h1ffb: x = 16'h25b1; 14'h1ffc: x = 16'h25b0; 14'h1ffd: x = 16'h25af; 14'h1ffe: x = 16'h25af; 14'h1fff: x = 16'h25ae; 14'h2000: x = 16'h25ad; 14'h2001: x = 16'h25ac; 14'h2002: x = 16'h25ab; 14'h2003: x = 16'h25aa; 14'h2004: x = 16'h25a9; 14'h2005: x = 16'h25a9; 14'h2006: x = 16'h25a8; 14'h2007: x = 16'h25a7; 14'h2008: x = 16'h25a6; 14'h2009: x = 16'h25a5; 14'h200a: x = 16'h25a4; 14'h200b: x = 16'h25a4; 14'h200c: x = 16'h25a3; 14'h200d: x = 16'h25a2; 14'h200e: x = 16'h25a1; 14'h200f: x = 16'h25a0; 14'h2010: x = 16'h259f; 14'h2011: x = 16'h259e; 14'h2012: x = 16'h259e; 14'h2013: x = 16'h259d; 14'h2014: x = 16'h259c; 14'h2015: x = 16'h259b; 14'h2016: x = 16'h259a; 14'h2017: x = 16'h2599; 14'h2018: x = 16'h2598; 14'h2019: x = 16'h2598; 14'h201a: x = 16'h2597; 14'h201b: x = 16'h2596; 14'h201c: x = 16'h2595; 14'h201d: x = 16'h2594; 14'h201e: x = 16'h2593; 14'h201f: x = 16'h2593; 14'h2020: x = 16'h2592; 14'h2021: x = 16'h2591; 14'h2022: x = 16'h2590; 14'h2023: x = 16'h258f; 14'h2024: x = 16'h258e; 14'h2025: x = 16'h258d; 14'h2026: x = 16'h258d; 14'h2027: x = 16'h258c; 14'h2028: x = 16'h258b; 14'h2029: x = 16'h258a; 14'h202a: x = 16'h2589; 14'h202b: x = 16'h2588; 14'h202c: x = 16'h2588; 14'h202d: x = 16'h2587; 14'h202e: x = 16'h2586; 14'h202f: x = 16'h2585; 14'h2030: x = 16'h2584; 14'h2031: x = 16'h2583; 14'h2032: x = 16'h2582; 14'h2033: x = 16'h2582; 14'h2034: x = 16'h2581; 14'h2035: x = 16'h2580; 14'h2036: x = 16'h257f; 14'h2037: x = 16'h257e; 14'h2038: x = 16'h257d; 14'h2039: x = 16'h257c; 14'h203a: x = 16'h257c; 14'h203b: x = 16'h257b; 14'h203c: x = 16'h257a; 14'h203d: x = 16'h2579; 14'h203e: x = 16'h2578; 14'h203f: x = 16'h2577; 14'h2040: x = 16'h2577; 14'h2041: x = 16'h2576; 14'h2042: x = 16'h2575; 14'h2043: x = 16'h2574; 14'h2044: x = 16'h2573; 14'h2045: x = 16'h2572; 14'h2046: x = 16'h2571; 14'h2047: x = 16'h2571; 14'h2048: x = 16'h2570; 14'h2049: x = 16'h256f; 14'h204a: x = 16'h256e; 14'h204b: x = 16'h256d; 14'h204c: x = 16'h256c; 14'h204d: x = 16'h256c; 14'h204e: x = 16'h256b; 14'h204f: x = 16'h256a; 14'h2050: x = 16'h2569; 14'h2051: x = 16'h2568; 14'h2052: x = 16'h2567; 14'h2053: x = 16'h2566; 14'h2054: x = 16'h2566; 14'h2055: x = 16'h2565; 14'h2056: x = 16'h2564; 14'h2057: x = 16'h2563; 14'h2058: x = 16'h2562; 14'h2059: x = 16'h2561; 14'h205a: x = 16'h2561; 14'h205b: x = 16'h2560; 14'h205c: x = 16'h255f; 14'h205d: x = 16'h255e; 14'h205e: x = 16'h255d; 14'h205f: x = 16'h255c; 14'h2060: x = 16'h255b; 14'h2061: x = 16'h255b; 14'h2062: x = 16'h255a; 14'h2063: x = 16'h2559; 14'h2064: x = 16'h2558; 14'h2065: x = 16'h2557; 14'h2066: x = 16'h2556; 14'h2067: x = 16'h2556; 14'h2068: x = 16'h2555; 14'h2069: x = 16'h2554; 14'h206a: x = 16'h2553; 14'h206b: x = 16'h2552; 14'h206c: x = 16'h2551; 14'h206d: x = 16'h2550; 14'h206e: x = 16'h2550; 14'h206f: x = 16'h254f; 14'h2070: x = 16'h254e; 14'h2071: x = 16'h254d; 14'h2072: x = 16'h254c; 14'h2073: x = 16'h254b; 14'h2074: x = 16'h254b; 14'h2075: x = 16'h254a; 14'h2076: x = 16'h2549; 14'h2077: x = 16'h2548; 14'h2078: x = 16'h2547; 14'h2079: x = 16'h2546; 14'h207a: x = 16'h2545; 14'h207b: x = 16'h2545; 14'h207c: x = 16'h2544; 14'h207d: x = 16'h2543; 14'h207e: x = 16'h2542; 14'h207f: x = 16'h2541; 14'h2080: x = 16'h2540; 14'h2081: x = 16'h2540; 14'h2082: x = 16'h253f; 14'h2083: x = 16'h253e; 14'h2084: x = 16'h253d; 14'h2085: x = 16'h253c; 14'h2086: x = 16'h253b; 14'h2087: x = 16'h253a; 14'h2088: x = 16'h253a; 14'h2089: x = 16'h2539; 14'h208a: x = 16'h2538; 14'h208b: x = 16'h2537; 14'h208c: x = 16'h2536; 14'h208d: x = 16'h2535; 14'h208e: x = 16'h2535; 14'h208f: x = 16'h2534; 14'h2090: x = 16'h2533; 14'h2091: x = 16'h2532; 14'h2092: x = 16'h2531; 14'h2093: x = 16'h2530; 14'h2094: x = 16'h252f; 14'h2095: x = 16'h252f; 14'h2096: x = 16'h252e; 14'h2097: x = 16'h252d; 14'h2098: x = 16'h252c; 14'h2099: x = 16'h252b; 14'h209a: x = 16'h252a; 14'h209b: x = 16'h252a; 14'h209c: x = 16'h2529; 14'h209d: x = 16'h2528; 14'h209e: x = 16'h2527; 14'h209f: x = 16'h2526; 14'h20a0: x = 16'h2525; 14'h20a1: x = 16'h2524; 14'h20a2: x = 16'h2524; 14'h20a3: x = 16'h2523; 14'h20a4: x = 16'h2522; 14'h20a5: x = 16'h2521; 14'h20a6: x = 16'h2520; 14'h20a7: x = 16'h251f; 14'h20a8: x = 16'h251f; 14'h20a9: x = 16'h251e; 14'h20aa: x = 16'h251d; 14'h20ab: x = 16'h251c; 14'h20ac: x = 16'h251b; 14'h20ad: x = 16'h251a; 14'h20ae: x = 16'h2519; 14'h20af: x = 16'h2519; 14'h20b0: x = 16'h2518; 14'h20b1: x = 16'h2517; 14'h20b2: x = 16'h2516; 14'h20b3: x = 16'h2515; 14'h20b4: x = 16'h2514; 14'h20b5: x = 16'h2514; 14'h20b6: x = 16'h2513; 14'h20b7: x = 16'h2512; 14'h20b8: x = 16'h2511; 14'h20b9: x = 16'h2510; 14'h20ba: x = 16'h250f; 14'h20bb: x = 16'h250f; 14'h20bc: x = 16'h250e; 14'h20bd: x = 16'h250d; 14'h20be: x = 16'h250c; 14'h20bf: x = 16'h250b; 14'h20c0: x = 16'h250a; 14'h20c1: x = 16'h2509; 14'h20c2: x = 16'h2509; 14'h20c3: x = 16'h2508; 14'h20c4: x = 16'h2507; 14'h20c5: x = 16'h2506; 14'h20c6: x = 16'h2505; 14'h20c7: x = 16'h2504; 14'h20c8: x = 16'h2504; 14'h20c9: x = 16'h2503; 14'h20ca: x = 16'h2502; 14'h20cb: x = 16'h2501; 14'h20cc: x = 16'h2500; 14'h20cd: x = 16'h24ff; 14'h20ce: x = 16'h24fe; 14'h20cf: x = 16'h24fe; 14'h20d0: x = 16'h24fd; 14'h20d1: x = 16'h24fc; 14'h20d2: x = 16'h24fb; 14'h20d3: x = 16'h24fa; 14'h20d4: x = 16'h24f9; 14'h20d5: x = 16'h24f9; 14'h20d6: x = 16'h24f8; 14'h20d7: x = 16'h24f7; 14'h20d8: x = 16'h24f6; 14'h20d9: x = 16'h24f5; 14'h20da: x = 16'h24f4; 14'h20db: x = 16'h24f4; 14'h20dc: x = 16'h24f3; 14'h20dd: x = 16'h24f2; 14'h20de: x = 16'h24f1; 14'h20df: x = 16'h24f0; 14'h20e0: x = 16'h24ef; 14'h20e1: x = 16'h24ee; 14'h20e2: x = 16'h24ee; 14'h20e3: x = 16'h24ed; 14'h20e4: x = 16'h24ec; 14'h20e5: x = 16'h24eb; 14'h20e6: x = 16'h24ea; 14'h20e7: x = 16'h24e9; 14'h20e8: x = 16'h24e9; 14'h20e9: x = 16'h24e8; 14'h20ea: x = 16'h24e7; 14'h20eb: x = 16'h24e6; 14'h20ec: x = 16'h24e5; 14'h20ed: x = 16'h24e4; 14'h20ee: x = 16'h24e3; 14'h20ef: x = 16'h24e3; 14'h20f0: x = 16'h24e2; 14'h20f1: x = 16'h24e1; 14'h20f2: x = 16'h24e0; 14'h20f3: x = 16'h24df; 14'h20f4: x = 16'h24de; 14'h20f5: x = 16'h24de; 14'h20f6: x = 16'h24dd; 14'h20f7: x = 16'h24dc; 14'h20f8: x = 16'h24db; 14'h20f9: x = 16'h24da; 14'h20fa: x = 16'h24d9; 14'h20fb: x = 16'h24d9; 14'h20fc: x = 16'h24d8; 14'h20fd: x = 16'h24d7; 14'h20fe: x = 16'h24d6; 14'h20ff: x = 16'h24d5; 14'h2100: x = 16'h24d4; 14'h2101: x = 16'h24d3; 14'h2102: x = 16'h24d3; 14'h2103: x = 16'h24d2; 14'h2104: x = 16'h24d1; 14'h2105: x = 16'h24d0; 14'h2106: x = 16'h24cf; 14'h2107: x = 16'h24ce; 14'h2108: x = 16'h24ce; 14'h2109: x = 16'h24cd; 14'h210a: x = 16'h24cc; 14'h210b: x = 16'h24cb; 14'h210c: x = 16'h24ca; 14'h210d: x = 16'h24c9; 14'h210e: x = 16'h24c9; 14'h210f: x = 16'h24c8; 14'h2110: x = 16'h24c7; 14'h2111: x = 16'h24c6; 14'h2112: x = 16'h24c5; 14'h2113: x = 16'h24c4; 14'h2114: x = 16'h24c3; 14'h2115: x = 16'h24c3; 14'h2116: x = 16'h24c2; 14'h2117: x = 16'h24c1; 14'h2118: x = 16'h24c0; 14'h2119: x = 16'h24bf; 14'h211a: x = 16'h24be; 14'h211b: x = 16'h24be; 14'h211c: x = 16'h24bd; 14'h211d: x = 16'h24bc; 14'h211e: x = 16'h24bb; 14'h211f: x = 16'h24ba; 14'h2120: x = 16'h24b9; 14'h2121: x = 16'h24b9; 14'h2122: x = 16'h24b8; 14'h2123: x = 16'h24b7; 14'h2124: x = 16'h24b6; 14'h2125: x = 16'h24b5; 14'h2126: x = 16'h24b4; 14'h2127: x = 16'h24b3; 14'h2128: x = 16'h24b3; 14'h2129: x = 16'h24b2; 14'h212a: x = 16'h24b1; 14'h212b: x = 16'h24b0; 14'h212c: x = 16'h24af; 14'h212d: x = 16'h24ae; 14'h212e: x = 16'h24ae; 14'h212f: x = 16'h24ad; 14'h2130: x = 16'h24ac; 14'h2131: x = 16'h24ab; 14'h2132: x = 16'h24aa; 14'h2133: x = 16'h24a9; 14'h2134: x = 16'h24a9; 14'h2135: x = 16'h24a8; 14'h2136: x = 16'h24a7; 14'h2137: x = 16'h24a6; 14'h2138: x = 16'h24a5; 14'h2139: x = 16'h24a4; 14'h213a: x = 16'h24a3; 14'h213b: x = 16'h24a3; 14'h213c: x = 16'h24a2; 14'h213d: x = 16'h24a1; 14'h213e: x = 16'h24a0; 14'h213f: x = 16'h249f; 14'h2140: x = 16'h249e; 14'h2141: x = 16'h249e; 14'h2142: x = 16'h249d; 14'h2143: x = 16'h249c; 14'h2144: x = 16'h249b; 14'h2145: x = 16'h249a; 14'h2146: x = 16'h2499; 14'h2147: x = 16'h2499; 14'h2148: x = 16'h2498; 14'h2149: x = 16'h2497; 14'h214a: x = 16'h2496; 14'h214b: x = 16'h2495; 14'h214c: x = 16'h2494; 14'h214d: x = 16'h2494; 14'h214e: x = 16'h2493; 14'h214f: x = 16'h2492; 14'h2150: x = 16'h2491; 14'h2151: x = 16'h2490; 14'h2152: x = 16'h248f; 14'h2153: x = 16'h248e; 14'h2154: x = 16'h248e; 14'h2155: x = 16'h248d; 14'h2156: x = 16'h248c; 14'h2157: x = 16'h248b; 14'h2158: x = 16'h248a; 14'h2159: x = 16'h2489; 14'h215a: x = 16'h2489; 14'h215b: x = 16'h2488; 14'h215c: x = 16'h2487; 14'h215d: x = 16'h2486; 14'h215e: x = 16'h2485; 14'h215f: x = 16'h2484; 14'h2160: x = 16'h2484; 14'h2161: x = 16'h2483; 14'h2162: x = 16'h2482; 14'h2163: x = 16'h2481; 14'h2164: x = 16'h2480; 14'h2165: x = 16'h247f; 14'h2166: x = 16'h247f; 14'h2167: x = 16'h247e; 14'h2168: x = 16'h247d; 14'h2169: x = 16'h247c; 14'h216a: x = 16'h247b; 14'h216b: x = 16'h247a; 14'h216c: x = 16'h2479; 14'h216d: x = 16'h2479; 14'h216e: x = 16'h2478; 14'h216f: x = 16'h2477; 14'h2170: x = 16'h2476; 14'h2171: x = 16'h2475; 14'h2172: x = 16'h2474; 14'h2173: x = 16'h2474; 14'h2174: x = 16'h2473; 14'h2175: x = 16'h2472; 14'h2176: x = 16'h2471; 14'h2177: x = 16'h2470; 14'h2178: x = 16'h246f; 14'h2179: x = 16'h246f; 14'h217a: x = 16'h246e; 14'h217b: x = 16'h246d; 14'h217c: x = 16'h246c; 14'h217d: x = 16'h246b; 14'h217e: x = 16'h246a; 14'h217f: x = 16'h246a; 14'h2180: x = 16'h2469; 14'h2181: x = 16'h2468; 14'h2182: x = 16'h2467; 14'h2183: x = 16'h2466; 14'h2184: x = 16'h2465; 14'h2185: x = 16'h2464; 14'h2186: x = 16'h2464; 14'h2187: x = 16'h2463; 14'h2188: x = 16'h2462; 14'h2189: x = 16'h2461; 14'h218a: x = 16'h2460; 14'h218b: x = 16'h245f; 14'h218c: x = 16'h245f; 14'h218d: x = 16'h245e; 14'h218e: x = 16'h245d; 14'h218f: x = 16'h245c; 14'h2190: x = 16'h245b; 14'h2191: x = 16'h245a; 14'h2192: x = 16'h245a; 14'h2193: x = 16'h2459; 14'h2194: x = 16'h2458; 14'h2195: x = 16'h2457; 14'h2196: x = 16'h2456; 14'h2197: x = 16'h2455; 14'h2198: x = 16'h2455; 14'h2199: x = 16'h2454; 14'h219a: x = 16'h2453; 14'h219b: x = 16'h2452; 14'h219c: x = 16'h2451; 14'h219d: x = 16'h2450; 14'h219e: x = 16'h244f; 14'h219f: x = 16'h244f; 14'h21a0: x = 16'h244e; 14'h21a1: x = 16'h244d; 14'h21a2: x = 16'h244c; 14'h21a3: x = 16'h244b; 14'h21a4: x = 16'h244a; 14'h21a5: x = 16'h244a; 14'h21a6: x = 16'h2449; 14'h21a7: x = 16'h2448; 14'h21a8: x = 16'h2447; 14'h21a9: x = 16'h2446; 14'h21aa: x = 16'h2445; 14'h21ab: x = 16'h2445; 14'h21ac: x = 16'h2444; 14'h21ad: x = 16'h2443; 14'h21ae: x = 16'h2442; 14'h21af: x = 16'h2441; 14'h21b0: x = 16'h2440; 14'h21b1: x = 16'h2440; 14'h21b2: x = 16'h243f; 14'h21b3: x = 16'h243e; 14'h21b4: x = 16'h243d; 14'h21b5: x = 16'h243c; 14'h21b6: x = 16'h243b; 14'h21b7: x = 16'h243b; 14'h21b8: x = 16'h243a; 14'h21b9: x = 16'h2439; 14'h21ba: x = 16'h2438; 14'h21bb: x = 16'h2437; 14'h21bc: x = 16'h2436; 14'h21bd: x = 16'h2435; 14'h21be: x = 16'h2435; 14'h21bf: x = 16'h2434; 14'h21c0: x = 16'h2433; 14'h21c1: x = 16'h2432; 14'h21c2: x = 16'h2431; 14'h21c3: x = 16'h2430; 14'h21c4: x = 16'h2430; 14'h21c5: x = 16'h242f; 14'h21c6: x = 16'h242e; 14'h21c7: x = 16'h242d; 14'h21c8: x = 16'h242c; 14'h21c9: x = 16'h242b; 14'h21ca: x = 16'h242b; 14'h21cb: x = 16'h242a; 14'h21cc: x = 16'h2429; 14'h21cd: x = 16'h2428; 14'h21ce: x = 16'h2427; 14'h21cf: x = 16'h2426; 14'h21d0: x = 16'h2426; 14'h21d1: x = 16'h2425; 14'h21d2: x = 16'h2424; 14'h21d3: x = 16'h2423; 14'h21d4: x = 16'h2422; 14'h21d5: x = 16'h2421; 14'h21d6: x = 16'h2421; 14'h21d7: x = 16'h2420; 14'h21d8: x = 16'h241f; 14'h21d9: x = 16'h241e; 14'h21da: x = 16'h241d; 14'h21db: x = 16'h241c; 14'h21dc: x = 16'h241c; 14'h21dd: x = 16'h241b; 14'h21de: x = 16'h241a; 14'h21df: x = 16'h2419; 14'h21e0: x = 16'h2418; 14'h21e1: x = 16'h2417; 14'h21e2: x = 16'h2417; 14'h21e3: x = 16'h2416; 14'h21e4: x = 16'h2415; 14'h21e5: x = 16'h2414; 14'h21e6: x = 16'h2413; 14'h21e7: x = 16'h2412; 14'h21e8: x = 16'h2411; 14'h21e9: x = 16'h2411; 14'h21ea: x = 16'h2410; 14'h21eb: x = 16'h240f; 14'h21ec: x = 16'h240e; 14'h21ed: x = 16'h240d; 14'h21ee: x = 16'h240c; 14'h21ef: x = 16'h240c; 14'h21f0: x = 16'h240b; 14'h21f1: x = 16'h240a; 14'h21f2: x = 16'h2409; 14'h21f3: x = 16'h2408; 14'h21f4: x = 16'h2407; 14'h21f5: x = 16'h2407; 14'h21f6: x = 16'h2406; 14'h21f7: x = 16'h2405; 14'h21f8: x = 16'h2404; 14'h21f9: x = 16'h2403; 14'h21fa: x = 16'h2402; 14'h21fb: x = 16'h2402; 14'h21fc: x = 16'h2401; 14'h21fd: x = 16'h2400; 14'h21fe: x = 16'h23ff; 14'h21ff: x = 16'h23fe; 14'h2200: x = 16'h23fd; 14'h2201: x = 16'h23fd; 14'h2202: x = 16'h23fc; 14'h2203: x = 16'h23fb; 14'h2204: x = 16'h23fa; 14'h2205: x = 16'h23f9; 14'h2206: x = 16'h23f8; 14'h2207: x = 16'h23f8; 14'h2208: x = 16'h23f7; 14'h2209: x = 16'h23f6; 14'h220a: x = 16'h23f5; 14'h220b: x = 16'h23f4; 14'h220c: x = 16'h23f3; 14'h220d: x = 16'h23f3; 14'h220e: x = 16'h23f2; 14'h220f: x = 16'h23f1; 14'h2210: x = 16'h23f0; 14'h2211: x = 16'h23ef; 14'h2212: x = 16'h23ee; 14'h2213: x = 16'h23ed; 14'h2214: x = 16'h23ed; 14'h2215: x = 16'h23ec; 14'h2216: x = 16'h23eb; 14'h2217: x = 16'h23ea; 14'h2218: x = 16'h23e9; 14'h2219: x = 16'h23e8; 14'h221a: x = 16'h23e8; 14'h221b: x = 16'h23e7; 14'h221c: x = 16'h23e6; 14'h221d: x = 16'h23e5; 14'h221e: x = 16'h23e4; 14'h221f: x = 16'h23e3; 14'h2220: x = 16'h23e3; 14'h2221: x = 16'h23e2; 14'h2222: x = 16'h23e1; 14'h2223: x = 16'h23e0; 14'h2224: x = 16'h23df; 14'h2225: x = 16'h23de; 14'h2226: x = 16'h23de; 14'h2227: x = 16'h23dd; 14'h2228: x = 16'h23dc; 14'h2229: x = 16'h23db; 14'h222a: x = 16'h23da; 14'h222b: x = 16'h23d9; 14'h222c: x = 16'h23d9; 14'h222d: x = 16'h23d8; 14'h222e: x = 16'h23d7; 14'h222f: x = 16'h23d6; 14'h2230: x = 16'h23d5; 14'h2231: x = 16'h23d4; 14'h2232: x = 16'h23d4; 14'h2233: x = 16'h23d3; 14'h2234: x = 16'h23d2; 14'h2235: x = 16'h23d1; 14'h2236: x = 16'h23d0; 14'h2237: x = 16'h23cf; 14'h2238: x = 16'h23cf; 14'h2239: x = 16'h23ce; 14'h223a: x = 16'h23cd; 14'h223b: x = 16'h23cc; 14'h223c: x = 16'h23cb; 14'h223d: x = 16'h23ca; 14'h223e: x = 16'h23ca; 14'h223f: x = 16'h23c9; 14'h2240: x = 16'h23c8; 14'h2241: x = 16'h23c7; 14'h2242: x = 16'h23c6; 14'h2243: x = 16'h23c5; 14'h2244: x = 16'h23c5; 14'h2245: x = 16'h23c4; 14'h2246: x = 16'h23c3; 14'h2247: x = 16'h23c2; 14'h2248: x = 16'h23c1; 14'h2249: x = 16'h23c0; 14'h224a: x = 16'h23c0; 14'h224b: x = 16'h23bf; 14'h224c: x = 16'h23be; 14'h224d: x = 16'h23bd; 14'h224e: x = 16'h23bc; 14'h224f: x = 16'h23bb; 14'h2250: x = 16'h23bb; 14'h2251: x = 16'h23ba; 14'h2252: x = 16'h23b9; 14'h2253: x = 16'h23b8; 14'h2254: x = 16'h23b7; 14'h2255: x = 16'h23b6; 14'h2256: x = 16'h23b5; 14'h2257: x = 16'h23b5; 14'h2258: x = 16'h23b4; 14'h2259: x = 16'h23b3; 14'h225a: x = 16'h23b2; 14'h225b: x = 16'h23b1; 14'h225c: x = 16'h23b0; 14'h225d: x = 16'h23b0; 14'h225e: x = 16'h23af; 14'h225f: x = 16'h23ae; 14'h2260: x = 16'h23ad; 14'h2261: x = 16'h23ac; 14'h2262: x = 16'h23ab; 14'h2263: x = 16'h23ab; 14'h2264: x = 16'h23aa; 14'h2265: x = 16'h23a9; 14'h2266: x = 16'h23a8; 14'h2267: x = 16'h23a7; 14'h2268: x = 16'h23a6; 14'h2269: x = 16'h23a6; 14'h226a: x = 16'h23a5; 14'h226b: x = 16'h23a4; 14'h226c: x = 16'h23a3; 14'h226d: x = 16'h23a2; 14'h226e: x = 16'h23a1; 14'h226f: x = 16'h23a1; 14'h2270: x = 16'h23a0; 14'h2271: x = 16'h239f; 14'h2272: x = 16'h239e; 14'h2273: x = 16'h239d; 14'h2274: x = 16'h239c; 14'h2275: x = 16'h239c; 14'h2276: x = 16'h239b; 14'h2277: x = 16'h239a; 14'h2278: x = 16'h2399; 14'h2279: x = 16'h2398; 14'h227a: x = 16'h2397; 14'h227b: x = 16'h2397; 14'h227c: x = 16'h2396; 14'h227d: x = 16'h2395; 14'h227e: x = 16'h2394; 14'h227f: x = 16'h2393; 14'h2280: x = 16'h2392; 14'h2281: x = 16'h2392; 14'h2282: x = 16'h2391; 14'h2283: x = 16'h2390; 14'h2284: x = 16'h238f; 14'h2285: x = 16'h238e; 14'h2286: x = 16'h238d; 14'h2287: x = 16'h238d; 14'h2288: x = 16'h238c; 14'h2289: x = 16'h238b; 14'h228a: x = 16'h238a; 14'h228b: x = 16'h2389; 14'h228c: x = 16'h2388; 14'h228d: x = 16'h2388; 14'h228e: x = 16'h2387; 14'h228f: x = 16'h2386; 14'h2290: x = 16'h2385; 14'h2291: x = 16'h2384; 14'h2292: x = 16'h2383; 14'h2293: x = 16'h2383; 14'h2294: x = 16'h2382; 14'h2295: x = 16'h2381; 14'h2296: x = 16'h2380; 14'h2297: x = 16'h237f; 14'h2298: x = 16'h237e; 14'h2299: x = 16'h237e; 14'h229a: x = 16'h237d; 14'h229b: x = 16'h237c; 14'h229c: x = 16'h237b; 14'h229d: x = 16'h237a; 14'h229e: x = 16'h2379; 14'h229f: x = 16'h2379; 14'h22a0: x = 16'h2378; 14'h22a1: x = 16'h2377; 14'h22a2: x = 16'h2376; 14'h22a3: x = 16'h2375; 14'h22a4: x = 16'h2374; 14'h22a5: x = 16'h2374; 14'h22a6: x = 16'h2373; 14'h22a7: x = 16'h2372; 14'h22a8: x = 16'h2371; 14'h22a9: x = 16'h2370; 14'h22aa: x = 16'h236f; 14'h22ab: x = 16'h236f; 14'h22ac: x = 16'h236e; 14'h22ad: x = 16'h236d; 14'h22ae: x = 16'h236c; 14'h22af: x = 16'h236b; 14'h22b0: x = 16'h236a; 14'h22b1: x = 16'h236a; 14'h22b2: x = 16'h2369; 14'h22b3: x = 16'h2368; 14'h22b4: x = 16'h2367; 14'h22b5: x = 16'h2366; 14'h22b6: x = 16'h2365; 14'h22b7: x = 16'h2365; 14'h22b8: x = 16'h2364; 14'h22b9: x = 16'h2363; 14'h22ba: x = 16'h2362; 14'h22bb: x = 16'h2361; 14'h22bc: x = 16'h2360; 14'h22bd: x = 16'h2360; 14'h22be: x = 16'h235f; 14'h22bf: x = 16'h235e; 14'h22c0: x = 16'h235d; 14'h22c1: x = 16'h235c; 14'h22c2: x = 16'h235b; 14'h22c3: x = 16'h235b; 14'h22c4: x = 16'h235a; 14'h22c5: x = 16'h2359; 14'h22c6: x = 16'h2358; 14'h22c7: x = 16'h2357; 14'h22c8: x = 16'h2356; 14'h22c9: x = 16'h2356; 14'h22ca: x = 16'h2355; 14'h22cb: x = 16'h2354; 14'h22cc: x = 16'h2353; 14'h22cd: x = 16'h2352; 14'h22ce: x = 16'h2351; 14'h22cf: x = 16'h2351; 14'h22d0: x = 16'h2350; 14'h22d1: x = 16'h234f; 14'h22d2: x = 16'h234e; 14'h22d3: x = 16'h234d; 14'h22d4: x = 16'h234c; 14'h22d5: x = 16'h234c; 14'h22d6: x = 16'h234b; 14'h22d7: x = 16'h234a; 14'h22d8: x = 16'h2349; 14'h22d9: x = 16'h2348; 14'h22da: x = 16'h2347; 14'h22db: x = 16'h2347; 14'h22dc: x = 16'h2346; 14'h22dd: x = 16'h2345; 14'h22de: x = 16'h2344; 14'h22df: x = 16'h2343; 14'h22e0: x = 16'h2342; 14'h22e1: x = 16'h2342; 14'h22e2: x = 16'h2341; 14'h22e3: x = 16'h2340; 14'h22e4: x = 16'h233f; 14'h22e5: x = 16'h233e; 14'h22e6: x = 16'h233d; 14'h22e7: x = 16'h233d; 14'h22e8: x = 16'h233c; 14'h22e9: x = 16'h233b; 14'h22ea: x = 16'h233a; 14'h22eb: x = 16'h2339; 14'h22ec: x = 16'h2338; 14'h22ed: x = 16'h2338; 14'h22ee: x = 16'h2337; 14'h22ef: x = 16'h2336; 14'h22f0: x = 16'h2335; 14'h22f1: x = 16'h2334; 14'h22f2: x = 16'h2333; 14'h22f3: x = 16'h2333; 14'h22f4: x = 16'h2332; 14'h22f5: x = 16'h2331; 14'h22f6: x = 16'h2330; 14'h22f7: x = 16'h232f; 14'h22f8: x = 16'h232e; 14'h22f9: x = 16'h232e; 14'h22fa: x = 16'h232d; 14'h22fb: x = 16'h232c; 14'h22fc: x = 16'h232b; 14'h22fd: x = 16'h232a; 14'h22fe: x = 16'h2329; 14'h22ff: x = 16'h2329; 14'h2300: x = 16'h2328; 14'h2301: x = 16'h2327; 14'h2302: x = 16'h2326; 14'h2303: x = 16'h2325; 14'h2304: x = 16'h2324; 14'h2305: x = 16'h2324; 14'h2306: x = 16'h2323; 14'h2307: x = 16'h2322; 14'h2308: x = 16'h2321; 14'h2309: x = 16'h2320; 14'h230a: x = 16'h231f; 14'h230b: x = 16'h231f; 14'h230c: x = 16'h231e; 14'h230d: x = 16'h231d; 14'h230e: x = 16'h231c; 14'h230f: x = 16'h231b; 14'h2310: x = 16'h231a; 14'h2311: x = 16'h231a; 14'h2312: x = 16'h2319; 14'h2313: x = 16'h2318; 14'h2314: x = 16'h2317; 14'h2315: x = 16'h2316; 14'h2316: x = 16'h2315; 14'h2317: x = 16'h2315; 14'h2318: x = 16'h2314; 14'h2319: x = 16'h2313; 14'h231a: x = 16'h2312; 14'h231b: x = 16'h2311; 14'h231c: x = 16'h2310; 14'h231d: x = 16'h2310; 14'h231e: x = 16'h230f; 14'h231f: x = 16'h230e; 14'h2320: x = 16'h230d; 14'h2321: x = 16'h230c; 14'h2322: x = 16'h230b; 14'h2323: x = 16'h230b; 14'h2324: x = 16'h230a; 14'h2325: x = 16'h2309; 14'h2326: x = 16'h2308; 14'h2327: x = 16'h2307; 14'h2328: x = 16'h2307; 14'h2329: x = 16'h2306; 14'h232a: x = 16'h2305; 14'h232b: x = 16'h2304; 14'h232c: x = 16'h2303; 14'h232d: x = 16'h2302; 14'h232e: x = 16'h2302; 14'h232f: x = 16'h2301; 14'h2330: x = 16'h2300; 14'h2331: x = 16'h22ff; 14'h2332: x = 16'h22fe; 14'h2333: x = 16'h22fd; 14'h2334: x = 16'h22fd; 14'h2335: x = 16'h22fc; 14'h2336: x = 16'h22fb; 14'h2337: x = 16'h22fa; 14'h2338: x = 16'h22f9; 14'h2339: x = 16'h22f8; 14'h233a: x = 16'h22f8; 14'h233b: x = 16'h22f7; 14'h233c: x = 16'h22f6; 14'h233d: x = 16'h22f5; 14'h233e: x = 16'h22f4; 14'h233f: x = 16'h22f3; 14'h2340: x = 16'h22f3; 14'h2341: x = 16'h22f2; 14'h2342: x = 16'h22f1; 14'h2343: x = 16'h22f0; 14'h2344: x = 16'h22ef; 14'h2345: x = 16'h22ee; 14'h2346: x = 16'h22ee; 14'h2347: x = 16'h22ed; 14'h2348: x = 16'h22ec; 14'h2349: x = 16'h22eb; 14'h234a: x = 16'h22ea; 14'h234b: x = 16'h22e9; 14'h234c: x = 16'h22e9; 14'h234d: x = 16'h22e8; 14'h234e: x = 16'h22e7; 14'h234f: x = 16'h22e6; 14'h2350: x = 16'h22e5; 14'h2351: x = 16'h22e4; 14'h2352: x = 16'h22e4; 14'h2353: x = 16'h22e3; 14'h2354: x = 16'h22e2; 14'h2355: x = 16'h22e1; 14'h2356: x = 16'h22e0; 14'h2357: x = 16'h22df; 14'h2358: x = 16'h22df; 14'h2359: x = 16'h22de; 14'h235a: x = 16'h22dd; 14'h235b: x = 16'h22dc; 14'h235c: x = 16'h22db; 14'h235d: x = 16'h22da; 14'h235e: x = 16'h22da; 14'h235f: x = 16'h22d9; 14'h2360: x = 16'h22d8; 14'h2361: x = 16'h22d7; 14'h2362: x = 16'h22d6; 14'h2363: x = 16'h22d5; 14'h2364: x = 16'h22d5; 14'h2365: x = 16'h22d4; 14'h2366: x = 16'h22d3; 14'h2367: x = 16'h22d2; 14'h2368: x = 16'h22d1; 14'h2369: x = 16'h22d0; 14'h236a: x = 16'h22d0; 14'h236b: x = 16'h22cf; 14'h236c: x = 16'h22ce; 14'h236d: x = 16'h22cd; 14'h236e: x = 16'h22cc; 14'h236f: x = 16'h22cc; 14'h2370: x = 16'h22cb; 14'h2371: x = 16'h22ca; 14'h2372: x = 16'h22c9; 14'h2373: x = 16'h22c8; 14'h2374: x = 16'h22c7; 14'h2375: x = 16'h22c7; 14'h2376: x = 16'h22c6; 14'h2377: x = 16'h22c5; 14'h2378: x = 16'h22c4; 14'h2379: x = 16'h22c3; 14'h237a: x = 16'h22c2; 14'h237b: x = 16'h22c2; 14'h237c: x = 16'h22c1; 14'h237d: x = 16'h22c0; 14'h237e: x = 16'h22bf; 14'h237f: x = 16'h22be; 14'h2380: x = 16'h22bd; 14'h2381: x = 16'h22bd; 14'h2382: x = 16'h22bc; 14'h2383: x = 16'h22bb; 14'h2384: x = 16'h22ba; 14'h2385: x = 16'h22b9; 14'h2386: x = 16'h22b8; 14'h2387: x = 16'h22b8; 14'h2388: x = 16'h22b7; 14'h2389: x = 16'h22b6; 14'h238a: x = 16'h22b5; 14'h238b: x = 16'h22b4; 14'h238c: x = 16'h22b3; 14'h238d: x = 16'h22b3; 14'h238e: x = 16'h22b2; 14'h238f: x = 16'h22b1; 14'h2390: x = 16'h22b0; 14'h2391: x = 16'h22af; 14'h2392: x = 16'h22ae; 14'h2393: x = 16'h22ae; 14'h2394: x = 16'h22ad; 14'h2395: x = 16'h22ac; 14'h2396: x = 16'h22ab; 14'h2397: x = 16'h22aa; 14'h2398: x = 16'h22a9; 14'h2399: x = 16'h22a9; 14'h239a: x = 16'h22a8; 14'h239b: x = 16'h22a7; 14'h239c: x = 16'h22a6; 14'h239d: x = 16'h22a5; 14'h239e: x = 16'h22a4; 14'h239f: x = 16'h22a4; 14'h23a0: x = 16'h22a3; 14'h23a1: x = 16'h22a2; 14'h23a2: x = 16'h22a1; 14'h23a3: x = 16'h22a0; 14'h23a4: x = 16'h22a0; 14'h23a5: x = 16'h229f; 14'h23a6: x = 16'h229e; 14'h23a7: x = 16'h229d; 14'h23a8: x = 16'h229c; 14'h23a9: x = 16'h229b; 14'h23aa: x = 16'h229b; 14'h23ab: x = 16'h229a; 14'h23ac: x = 16'h2299; 14'h23ad: x = 16'h2298; 14'h23ae: x = 16'h2297; 14'h23af: x = 16'h2296; 14'h23b0: x = 16'h2296; 14'h23b1: x = 16'h2295; 14'h23b2: x = 16'h2294; 14'h23b3: x = 16'h2293; 14'h23b4: x = 16'h2292; 14'h23b5: x = 16'h2291; 14'h23b6: x = 16'h2291; 14'h23b7: x = 16'h2290; 14'h23b8: x = 16'h228f; 14'h23b9: x = 16'h228e; 14'h23ba: x = 16'h228d; 14'h23bb: x = 16'h228c; 14'h23bc: x = 16'h228c; 14'h23bd: x = 16'h228b; 14'h23be: x = 16'h228a; 14'h23bf: x = 16'h2289; 14'h23c0: x = 16'h2288; 14'h23c1: x = 16'h2287; 14'h23c2: x = 16'h2287; 14'h23c3: x = 16'h2286; 14'h23c4: x = 16'h2285; 14'h23c5: x = 16'h2284; 14'h23c6: x = 16'h2283; 14'h23c7: x = 16'h2282; 14'h23c8: x = 16'h2282; 14'h23c9: x = 16'h2281; 14'h23ca: x = 16'h2280; 14'h23cb: x = 16'h227f; 14'h23cc: x = 16'h227e; 14'h23cd: x = 16'h227d; 14'h23ce: x = 16'h227d; 14'h23cf: x = 16'h227c; 14'h23d0: x = 16'h227b; 14'h23d1: x = 16'h227a; 14'h23d2: x = 16'h2279; 14'h23d3: x = 16'h2279; 14'h23d4: x = 16'h2278; 14'h23d5: x = 16'h2277; 14'h23d6: x = 16'h2276; 14'h23d7: x = 16'h2275; 14'h23d8: x = 16'h2274; 14'h23d9: x = 16'h2274; 14'h23da: x = 16'h2273; 14'h23db: x = 16'h2272; 14'h23dc: x = 16'h2271; 14'h23dd: x = 16'h2270; 14'h23de: x = 16'h226f; 14'h23df: x = 16'h226f; 14'h23e0: x = 16'h226e; 14'h23e1: x = 16'h226d; 14'h23e2: x = 16'h226c; 14'h23e3: x = 16'h226b; 14'h23e4: x = 16'h226a; 14'h23e5: x = 16'h226a; 14'h23e6: x = 16'h2269; 14'h23e7: x = 16'h2268; 14'h23e8: x = 16'h2267; 14'h23e9: x = 16'h2266; 14'h23ea: x = 16'h2265; 14'h23eb: x = 16'h2265; 14'h23ec: x = 16'h2264; 14'h23ed: x = 16'h2263; 14'h23ee: x = 16'h2262; 14'h23ef: x = 16'h2261; 14'h23f0: x = 16'h2260; 14'h23f1: x = 16'h2260; 14'h23f2: x = 16'h225f; 14'h23f3: x = 16'h225e; 14'h23f4: x = 16'h225d; 14'h23f5: x = 16'h225c; 14'h23f6: x = 16'h225c; 14'h23f7: x = 16'h225b; 14'h23f8: x = 16'h225a; 14'h23f9: x = 16'h2259; 14'h23fa: x = 16'h2258; 14'h23fb: x = 16'h2257; 14'h23fc: x = 16'h2257; 14'h23fd: x = 16'h2256; 14'h23fe: x = 16'h2255; 14'h23ff: x = 16'h2254; 14'h2400: x = 16'h2253; 14'h2401: x = 16'h2252; 14'h2402: x = 16'h2252; 14'h2403: x = 16'h2251; 14'h2404: x = 16'h2250; 14'h2405: x = 16'h224f; 14'h2406: x = 16'h224e; 14'h2407: x = 16'h224d; 14'h2408: x = 16'h224d; 14'h2409: x = 16'h224c; 14'h240a: x = 16'h224b; 14'h240b: x = 16'h224a; 14'h240c: x = 16'h2249; 14'h240d: x = 16'h2248; 14'h240e: x = 16'h2248; 14'h240f: x = 16'h2247; 14'h2410: x = 16'h2246; 14'h2411: x = 16'h2245; 14'h2412: x = 16'h2244; 14'h2413: x = 16'h2243; 14'h2414: x = 16'h2243; 14'h2415: x = 16'h2242; 14'h2416: x = 16'h2241; 14'h2417: x = 16'h2240; 14'h2418: x = 16'h223f; 14'h2419: x = 16'h223f; 14'h241a: x = 16'h223e; 14'h241b: x = 16'h223d; 14'h241c: x = 16'h223c; 14'h241d: x = 16'h223b; 14'h241e: x = 16'h223a; 14'h241f: x = 16'h223a; 14'h2420: x = 16'h2239; 14'h2421: x = 16'h2238; 14'h2422: x = 16'h2237; 14'h2423: x = 16'h2236; 14'h2424: x = 16'h2235; 14'h2425: x = 16'h2235; 14'h2426: x = 16'h2234; 14'h2427: x = 16'h2233; 14'h2428: x = 16'h2232; 14'h2429: x = 16'h2231; 14'h242a: x = 16'h2230; 14'h242b: x = 16'h2230; 14'h242c: x = 16'h222f; 14'h242d: x = 16'h222e; 14'h242e: x = 16'h222d; 14'h242f: x = 16'h222c; 14'h2430: x = 16'h222b; 14'h2431: x = 16'h222b; 14'h2432: x = 16'h222a; 14'h2433: x = 16'h2229; 14'h2434: x = 16'h2228; 14'h2435: x = 16'h2227; 14'h2436: x = 16'h2226; 14'h2437: x = 16'h2226; 14'h2438: x = 16'h2225; 14'h2439: x = 16'h2224; 14'h243a: x = 16'h2223; 14'h243b: x = 16'h2222; 14'h243c: x = 16'h2222; 14'h243d: x = 16'h2221; 14'h243e: x = 16'h2220; 14'h243f: x = 16'h221f; 14'h2440: x = 16'h221e; 14'h2441: x = 16'h221d; 14'h2442: x = 16'h221d; 14'h2443: x = 16'h221c; 14'h2444: x = 16'h221b; 14'h2445: x = 16'h221a; 14'h2446: x = 16'h2219; 14'h2447: x = 16'h2218; 14'h2448: x = 16'h2218; 14'h2449: x = 16'h2217; 14'h244a: x = 16'h2216; 14'h244b: x = 16'h2215; 14'h244c: x = 16'h2214; 14'h244d: x = 16'h2213; 14'h244e: x = 16'h2213; 14'h244f: x = 16'h2212; 14'h2450: x = 16'h2211; 14'h2451: x = 16'h2210; 14'h2452: x = 16'h220f; 14'h2453: x = 16'h220e; 14'h2454: x = 16'h220e; 14'h2455: x = 16'h220d; 14'h2456: x = 16'h220c; 14'h2457: x = 16'h220b; 14'h2458: x = 16'h220a; 14'h2459: x = 16'h220a; 14'h245a: x = 16'h2209; 14'h245b: x = 16'h2208; 14'h245c: x = 16'h2207; 14'h245d: x = 16'h2206; 14'h245e: x = 16'h2205; 14'h245f: x = 16'h2205; 14'h2460: x = 16'h2204; 14'h2461: x = 16'h2203; 14'h2462: x = 16'h2202; 14'h2463: x = 16'h2201; 14'h2464: x = 16'h2200; 14'h2465: x = 16'h2200; 14'h2466: x = 16'h21ff; 14'h2467: x = 16'h21fe; 14'h2468: x = 16'h21fd; 14'h2469: x = 16'h21fc; 14'h246a: x = 16'h21fb; 14'h246b: x = 16'h21fb; 14'h246c: x = 16'h21fa; 14'h246d: x = 16'h21f9; 14'h246e: x = 16'h21f8; 14'h246f: x = 16'h21f7; 14'h2470: x = 16'h21f6; 14'h2471: x = 16'h21f6; 14'h2472: x = 16'h21f5; 14'h2473: x = 16'h21f4; 14'h2474: x = 16'h21f3; 14'h2475: x = 16'h21f2; 14'h2476: x = 16'h21f2; 14'h2477: x = 16'h21f1; 14'h2478: x = 16'h21f0; 14'h2479: x = 16'h21ef; 14'h247a: x = 16'h21ee; 14'h247b: x = 16'h21ed; 14'h247c: x = 16'h21ed; 14'h247d: x = 16'h21ec; 14'h247e: x = 16'h21eb; 14'h247f: x = 16'h21ea; 14'h2480: x = 16'h21e9; 14'h2481: x = 16'h21e8; 14'h2482: x = 16'h21e8; 14'h2483: x = 16'h21e7; 14'h2484: x = 16'h21e6; 14'h2485: x = 16'h21e5; 14'h2486: x = 16'h21e4; 14'h2487: x = 16'h21e3; 14'h2488: x = 16'h21e3; 14'h2489: x = 16'h21e2; 14'h248a: x = 16'h21e1; 14'h248b: x = 16'h21e0; 14'h248c: x = 16'h21df; 14'h248d: x = 16'h21de; 14'h248e: x = 16'h21de; 14'h248f: x = 16'h21dd; 14'h2490: x = 16'h21dc; 14'h2491: x = 16'h21db; 14'h2492: x = 16'h21da; 14'h2493: x = 16'h21da; 14'h2494: x = 16'h21d9; 14'h2495: x = 16'h21d8; 14'h2496: x = 16'h21d7; 14'h2497: x = 16'h21d6; 14'h2498: x = 16'h21d5; 14'h2499: x = 16'h21d5; 14'h249a: x = 16'h21d4; 14'h249b: x = 16'h21d3; 14'h249c: x = 16'h21d2; 14'h249d: x = 16'h21d1; 14'h249e: x = 16'h21d0; 14'h249f: x = 16'h21d0; 14'h24a0: x = 16'h21cf; 14'h24a1: x = 16'h21ce; 14'h24a2: x = 16'h21cd; 14'h24a3: x = 16'h21cc; 14'h24a4: x = 16'h21cb; 14'h24a5: x = 16'h21cb; 14'h24a6: x = 16'h21ca; 14'h24a7: x = 16'h21c9; 14'h24a8: x = 16'h21c8; 14'h24a9: x = 16'h21c7; 14'h24aa: x = 16'h21c7; 14'h24ab: x = 16'h21c6; 14'h24ac: x = 16'h21c5; 14'h24ad: x = 16'h21c4; 14'h24ae: x = 16'h21c3; 14'h24af: x = 16'h21c2; 14'h24b0: x = 16'h21c2; 14'h24b1: x = 16'h21c1; 14'h24b2: x = 16'h21c0; 14'h24b3: x = 16'h21bf; 14'h24b4: x = 16'h21be; 14'h24b5: x = 16'h21bd; 14'h24b6: x = 16'h21bd; 14'h24b7: x = 16'h21bc; 14'h24b8: x = 16'h21bb; 14'h24b9: x = 16'h21ba; 14'h24ba: x = 16'h21b9; 14'h24bb: x = 16'h21b8; 14'h24bc: x = 16'h21b8; 14'h24bd: x = 16'h21b7; 14'h24be: x = 16'h21b6; 14'h24bf: x = 16'h21b5; 14'h24c0: x = 16'h21b4; 14'h24c1: x = 16'h21b3; 14'h24c2: x = 16'h21b3; 14'h24c3: x = 16'h21b2; 14'h24c4: x = 16'h21b1; 14'h24c5: x = 16'h21b0; 14'h24c6: x = 16'h21af; 14'h24c7: x = 16'h21af; 14'h24c8: x = 16'h21ae; 14'h24c9: x = 16'h21ad; 14'h24ca: x = 16'h21ac; 14'h24cb: x = 16'h21ab; 14'h24cc: x = 16'h21aa; 14'h24cd: x = 16'h21aa; 14'h24ce: x = 16'h21a9; 14'h24cf: x = 16'h21a8; 14'h24d0: x = 16'h21a7; 14'h24d1: x = 16'h21a6; 14'h24d2: x = 16'h21a5; 14'h24d3: x = 16'h21a5; 14'h24d4: x = 16'h21a4; 14'h24d5: x = 16'h21a3; 14'h24d6: x = 16'h21a2; 14'h24d7: x = 16'h21a1; 14'h24d8: x = 16'h21a0; 14'h24d9: x = 16'h21a0; 14'h24da: x = 16'h219f; 14'h24db: x = 16'h219e; 14'h24dc: x = 16'h219d; 14'h24dd: x = 16'h219c; 14'h24de: x = 16'h219c; 14'h24df: x = 16'h219b; 14'h24e0: x = 16'h219a; 14'h24e1: x = 16'h2199; 14'h24e2: x = 16'h2198; 14'h24e3: x = 16'h2197; 14'h24e4: x = 16'h2197; 14'h24e5: x = 16'h2196; 14'h24e6: x = 16'h2195; 14'h24e7: x = 16'h2194; 14'h24e8: x = 16'h2193; 14'h24e9: x = 16'h2192; 14'h24ea: x = 16'h2192; 14'h24eb: x = 16'h2191; 14'h24ec: x = 16'h2190; 14'h24ed: x = 16'h218f; 14'h24ee: x = 16'h218e; 14'h24ef: x = 16'h218d; 14'h24f0: x = 16'h218d; 14'h24f1: x = 16'h218c; 14'h24f2: x = 16'h218b; 14'h24f3: x = 16'h218a; 14'h24f4: x = 16'h2189; 14'h24f5: x = 16'h2189; 14'h24f6: x = 16'h2188; 14'h24f7: x = 16'h2187; 14'h24f8: x = 16'h2186; 14'h24f9: x = 16'h2185; 14'h24fa: x = 16'h2184; 14'h24fb: x = 16'h2184; 14'h24fc: x = 16'h2183; 14'h24fd: x = 16'h2182; 14'h24fe: x = 16'h2181; 14'h24ff: x = 16'h2180; 14'h2500: x = 16'h217f; 14'h2501: x = 16'h217f; 14'h2502: x = 16'h217e; 14'h2503: x = 16'h217d; 14'h2504: x = 16'h217c; 14'h2505: x = 16'h217b; 14'h2506: x = 16'h217a; 14'h2507: x = 16'h217a; 14'h2508: x = 16'h2179; 14'h2509: x = 16'h2178; 14'h250a: x = 16'h2177; 14'h250b: x = 16'h2176; 14'h250c: x = 16'h2176; 14'h250d: x = 16'h2175; 14'h250e: x = 16'h2174; 14'h250f: x = 16'h2173; 14'h2510: x = 16'h2172; 14'h2511: x = 16'h2171; 14'h2512: x = 16'h2171; 14'h2513: x = 16'h2170; 14'h2514: x = 16'h216f; 14'h2515: x = 16'h216e; 14'h2516: x = 16'h216d; 14'h2517: x = 16'h216c; 14'h2518: x = 16'h216c; 14'h2519: x = 16'h216b; 14'h251a: x = 16'h216a; 14'h251b: x = 16'h2169; 14'h251c: x = 16'h2168; 14'h251d: x = 16'h2167; 14'h251e: x = 16'h2167; 14'h251f: x = 16'h2166; 14'h2520: x = 16'h2165; 14'h2521: x = 16'h2164; 14'h2522: x = 16'h2163; 14'h2523: x = 16'h2163; 14'h2524: x = 16'h2162; 14'h2525: x = 16'h2161; 14'h2526: x = 16'h2160; 14'h2527: x = 16'h215f; 14'h2528: x = 16'h215e; 14'h2529: x = 16'h215e; 14'h252a: x = 16'h215d; 14'h252b: x = 16'h215c; 14'h252c: x = 16'h215b; 14'h252d: x = 16'h215a; 14'h252e: x = 16'h2159; 14'h252f: x = 16'h2159; 14'h2530: x = 16'h2158; 14'h2531: x = 16'h2157; 14'h2532: x = 16'h2156; 14'h2533: x = 16'h2155; 14'h2534: x = 16'h2154; 14'h2535: x = 16'h2154; 14'h2536: x = 16'h2153; 14'h2537: x = 16'h2152; 14'h2538: x = 16'h2151; 14'h2539: x = 16'h2150; 14'h253a: x = 16'h2150; 14'h253b: x = 16'h214f; 14'h253c: x = 16'h214e; 14'h253d: x = 16'h214d; 14'h253e: x = 16'h214c; 14'h253f: x = 16'h214b; 14'h2540: x = 16'h214b; 14'h2541: x = 16'h214a; 14'h2542: x = 16'h2149; 14'h2543: x = 16'h2148; 14'h2544: x = 16'h2147; 14'h2545: x = 16'h2146; 14'h2546: x = 16'h2146; 14'h2547: x = 16'h2145; 14'h2548: x = 16'h2144; 14'h2549: x = 16'h2143; 14'h254a: x = 16'h2142; 14'h254b: x = 16'h2141; 14'h254c: x = 16'h2141; 14'h254d: x = 16'h2140; 14'h254e: x = 16'h213f; 14'h254f: x = 16'h213e; 14'h2550: x = 16'h213d; 14'h2551: x = 16'h213d; 14'h2552: x = 16'h213c; 14'h2553: x = 16'h213b; 14'h2554: x = 16'h213a; 14'h2555: x = 16'h2139; 14'h2556: x = 16'h2138; 14'h2557: x = 16'h2138; 14'h2558: x = 16'h2137; 14'h2559: x = 16'h2136; 14'h255a: x = 16'h2135; 14'h255b: x = 16'h2134; 14'h255c: x = 16'h2133; 14'h255d: x = 16'h2133; 14'h255e: x = 16'h2132; 14'h255f: x = 16'h2131; 14'h2560: x = 16'h2130; 14'h2561: x = 16'h212f; 14'h2562: x = 16'h212f; 14'h2563: x = 16'h212e; 14'h2564: x = 16'h212d; 14'h2565: x = 16'h212c; 14'h2566: x = 16'h212b; 14'h2567: x = 16'h212a; 14'h2568: x = 16'h212a; 14'h2569: x = 16'h2129; 14'h256a: x = 16'h2128; 14'h256b: x = 16'h2127; 14'h256c: x = 16'h2126; 14'h256d: x = 16'h2125; 14'h256e: x = 16'h2125; 14'h256f: x = 16'h2124; 14'h2570: x = 16'h2123; 14'h2571: x = 16'h2122; 14'h2572: x = 16'h2121; 14'h2573: x = 16'h2120; 14'h2574: x = 16'h2120; 14'h2575: x = 16'h211f; 14'h2576: x = 16'h211e; 14'h2577: x = 16'h211d; 14'h2578: x = 16'h211c; 14'h2579: x = 16'h211c; 14'h257a: x = 16'h211b; 14'h257b: x = 16'h211a; 14'h257c: x = 16'h2119; 14'h257d: x = 16'h2118; 14'h257e: x = 16'h2117; 14'h257f: x = 16'h2117; 14'h2580: x = 16'h2116; 14'h2581: x = 16'h2115; 14'h2582: x = 16'h2114; 14'h2583: x = 16'h2113; 14'h2584: x = 16'h2112; 14'h2585: x = 16'h2112; 14'h2586: x = 16'h2111; 14'h2587: x = 16'h2110; 14'h2588: x = 16'h210f; 14'h2589: x = 16'h210e; 14'h258a: x = 16'h210d; 14'h258b: x = 16'h210d; 14'h258c: x = 16'h210c; 14'h258d: x = 16'h210b; 14'h258e: x = 16'h210a; 14'h258f: x = 16'h2109; 14'h2590: x = 16'h2109; 14'h2591: x = 16'h2108; 14'h2592: x = 16'h2107; 14'h2593: x = 16'h2106; 14'h2594: x = 16'h2105; 14'h2595: x = 16'h2104; 14'h2596: x = 16'h2104; 14'h2597: x = 16'h2103; 14'h2598: x = 16'h2102; 14'h2599: x = 16'h2101; 14'h259a: x = 16'h2100; 14'h259b: x = 16'h20ff; 14'h259c: x = 16'h20ff; 14'h259d: x = 16'h20fe; 14'h259e: x = 16'h20fd; 14'h259f: x = 16'h20fc; 14'h25a0: x = 16'h20fb; 14'h25a1: x = 16'h20fb; 14'h25a2: x = 16'h20fa; 14'h25a3: x = 16'h20f9; 14'h25a4: x = 16'h20f8; 14'h25a5: x = 16'h20f7; 14'h25a6: x = 16'h20f6; 14'h25a7: x = 16'h20f6; 14'h25a8: x = 16'h20f5; 14'h25a9: x = 16'h20f4; 14'h25aa: x = 16'h20f3; 14'h25ab: x = 16'h20f2; 14'h25ac: x = 16'h20f1; 14'h25ad: x = 16'h20f1; 14'h25ae: x = 16'h20f0; 14'h25af: x = 16'h20ef; 14'h25b0: x = 16'h20ee; 14'h25b1: x = 16'h20ed; 14'h25b2: x = 16'h20ec; 14'h25b3: x = 16'h20ec; 14'h25b4: x = 16'h20eb; 14'h25b5: x = 16'h20ea; 14'h25b6: x = 16'h20e9; 14'h25b7: x = 16'h20e8; 14'h25b8: x = 16'h20e8; 14'h25b9: x = 16'h20e7; 14'h25ba: x = 16'h20e6; 14'h25bb: x = 16'h20e5; 14'h25bc: x = 16'h20e4; 14'h25bd: x = 16'h20e3; 14'h25be: x = 16'h20e3; 14'h25bf: x = 16'h20e2; 14'h25c0: x = 16'h20e1; 14'h25c1: x = 16'h20e0; 14'h25c2: x = 16'h20df; 14'h25c3: x = 16'h20de; 14'h25c4: x = 16'h20de; 14'h25c5: x = 16'h20dd; 14'h25c6: x = 16'h20dc; 14'h25c7: x = 16'h20db; 14'h25c8: x = 16'h20da; 14'h25c9: x = 16'h20da; 14'h25ca: x = 16'h20d9; 14'h25cb: x = 16'h20d8; 14'h25cc: x = 16'h20d7; 14'h25cd: x = 16'h20d6; 14'h25ce: x = 16'h20d5; 14'h25cf: x = 16'h20d5; 14'h25d0: x = 16'h20d4; 14'h25d1: x = 16'h20d3; 14'h25d2: x = 16'h20d2; 14'h25d3: x = 16'h20d1; 14'h25d4: x = 16'h20d0; 14'h25d5: x = 16'h20d0; 14'h25d6: x = 16'h20cf; 14'h25d7: x = 16'h20ce; 14'h25d8: x = 16'h20cd; 14'h25d9: x = 16'h20cc; 14'h25da: x = 16'h20cb; 14'h25db: x = 16'h20cb; 14'h25dc: x = 16'h20ca; 14'h25dd: x = 16'h20c9; 14'h25de: x = 16'h20c8; 14'h25df: x = 16'h20c7; 14'h25e0: x = 16'h20c7; 14'h25e1: x = 16'h20c6; 14'h25e2: x = 16'h20c5; 14'h25e3: x = 16'h20c4; 14'h25e4: x = 16'h20c3; 14'h25e5: x = 16'h20c2; 14'h25e6: x = 16'h20c2; 14'h25e7: x = 16'h20c1; 14'h25e8: x = 16'h20c0; 14'h25e9: x = 16'h20bf; 14'h25ea: x = 16'h20be; 14'h25eb: x = 16'h20bd; 14'h25ec: x = 16'h20bd; 14'h25ed: x = 16'h20bc; 14'h25ee: x = 16'h20bb; 14'h25ef: x = 16'h20ba; 14'h25f0: x = 16'h20b9; 14'h25f1: x = 16'h20b9; 14'h25f2: x = 16'h20b8; 14'h25f3: x = 16'h20b7; 14'h25f4: x = 16'h20b6; 14'h25f5: x = 16'h20b5; 14'h25f6: x = 16'h20b4; 14'h25f7: x = 16'h20b4; 14'h25f8: x = 16'h20b3; 14'h25f9: x = 16'h20b2; 14'h25fa: x = 16'h20b1; 14'h25fb: x = 16'h20b0; 14'h25fc: x = 16'h20af; 14'h25fd: x = 16'h20af; 14'h25fe: x = 16'h20ae; 14'h25ff: x = 16'h20ad; 14'h2600: x = 16'h20ac; 14'h2601: x = 16'h20ab; 14'h2602: x = 16'h20aa; 14'h2603: x = 16'h20aa; 14'h2604: x = 16'h20a9; 14'h2605: x = 16'h20a8; 14'h2606: x = 16'h20a7; 14'h2607: x = 16'h20a6; 14'h2608: x = 16'h20a6; 14'h2609: x = 16'h20a5; 14'h260a: x = 16'h20a4; 14'h260b: x = 16'h20a3; 14'h260c: x = 16'h20a2; 14'h260d: x = 16'h20a1; 14'h260e: x = 16'h20a1; 14'h260f: x = 16'h20a0; 14'h2610: x = 16'h209f; 14'h2611: x = 16'h209e; 14'h2612: x = 16'h209d; 14'h2613: x = 16'h209c; 14'h2614: x = 16'h209c; 14'h2615: x = 16'h209b; 14'h2616: x = 16'h209a; 14'h2617: x = 16'h2099; 14'h2618: x = 16'h2098; 14'h2619: x = 16'h2098; 14'h261a: x = 16'h2097; 14'h261b: x = 16'h2096; 14'h261c: x = 16'h2095; 14'h261d: x = 16'h2094; 14'h261e: x = 16'h2093; 14'h261f: x = 16'h2093; 14'h2620: x = 16'h2092; 14'h2621: x = 16'h2091; 14'h2622: x = 16'h2090; 14'h2623: x = 16'h208f; 14'h2624: x = 16'h208e; 14'h2625: x = 16'h208e; 14'h2626: x = 16'h208d; 14'h2627: x = 16'h208c; 14'h2628: x = 16'h208b; 14'h2629: x = 16'h208a; 14'h262a: x = 16'h208a; 14'h262b: x = 16'h2089; 14'h262c: x = 16'h2088; 14'h262d: x = 16'h2087; 14'h262e: x = 16'h2086; 14'h262f: x = 16'h2085; 14'h2630: x = 16'h2085; 14'h2631: x = 16'h2084; 14'h2632: x = 16'h2083; 14'h2633: x = 16'h2082; 14'h2634: x = 16'h2081; 14'h2635: x = 16'h2080; 14'h2636: x = 16'h2080; 14'h2637: x = 16'h207f; 14'h2638: x = 16'h207e; 14'h2639: x = 16'h207d; 14'h263a: x = 16'h207c; 14'h263b: x = 16'h207b; 14'h263c: x = 16'h207b; 14'h263d: x = 16'h207a; 14'h263e: x = 16'h2079; 14'h263f: x = 16'h2078; 14'h2640: x = 16'h2077; 14'h2641: x = 16'h2077; 14'h2642: x = 16'h2076; 14'h2643: x = 16'h2075; 14'h2644: x = 16'h2074; 14'h2645: x = 16'h2073; 14'h2646: x = 16'h2072; 14'h2647: x = 16'h2072; 14'h2648: x = 16'h2071; 14'h2649: x = 16'h2070; 14'h264a: x = 16'h206f; 14'h264b: x = 16'h206e; 14'h264c: x = 16'h206d; 14'h264d: x = 16'h206d; 14'h264e: x = 16'h206c; 14'h264f: x = 16'h206b; 14'h2650: x = 16'h206a; 14'h2651: x = 16'h2069; 14'h2652: x = 16'h2069; 14'h2653: x = 16'h2068; 14'h2654: x = 16'h2067; 14'h2655: x = 16'h2066; 14'h2656: x = 16'h2065; 14'h2657: x = 16'h2064; 14'h2658: x = 16'h2064; 14'h2659: x = 16'h2063; 14'h265a: x = 16'h2062; 14'h265b: x = 16'h2061; 14'h265c: x = 16'h2060; 14'h265d: x = 16'h205f; 14'h265e: x = 16'h205f; 14'h265f: x = 16'h205e; 14'h2660: x = 16'h205d; 14'h2661: x = 16'h205c; 14'h2662: x = 16'h205b; 14'h2663: x = 16'h205b; 14'h2664: x = 16'h205a; 14'h2665: x = 16'h2059; 14'h2666: x = 16'h2058; 14'h2667: x = 16'h2057; 14'h2668: x = 16'h2056; 14'h2669: x = 16'h2056; 14'h266a: x = 16'h2055; 14'h266b: x = 16'h2054; 14'h266c: x = 16'h2053; 14'h266d: x = 16'h2052; 14'h266e: x = 16'h2051; 14'h266f: x = 16'h2051; 14'h2670: x = 16'h2050; 14'h2671: x = 16'h204f; 14'h2672: x = 16'h204e; 14'h2673: x = 16'h204d; 14'h2674: x = 16'h204c; 14'h2675: x = 16'h204c; 14'h2676: x = 16'h204b; 14'h2677: x = 16'h204a; 14'h2678: x = 16'h2049; 14'h2679: x = 16'h2048; 14'h267a: x = 16'h2048; 14'h267b: x = 16'h2047; 14'h267c: x = 16'h2046; 14'h267d: x = 16'h2045; 14'h267e: x = 16'h2044; 14'h267f: x = 16'h2043; 14'h2680: x = 16'h2043; 14'h2681: x = 16'h2042; 14'h2682: x = 16'h2041; 14'h2683: x = 16'h2040; 14'h2684: x = 16'h203f; 14'h2685: x = 16'h203e; 14'h2686: x = 16'h203e; 14'h2687: x = 16'h203d; 14'h2688: x = 16'h203c; 14'h2689: x = 16'h203b; 14'h268a: x = 16'h203a; 14'h268b: x = 16'h203a; 14'h268c: x = 16'h2039; 14'h268d: x = 16'h2038; 14'h268e: x = 16'h2037; 14'h268f: x = 16'h2036; 14'h2690: x = 16'h2035; 14'h2691: x = 16'h2035; 14'h2692: x = 16'h2034; 14'h2693: x = 16'h2033; 14'h2694: x = 16'h2032; 14'h2695: x = 16'h2031; 14'h2696: x = 16'h2030; 14'h2697: x = 16'h2030; 14'h2698: x = 16'h202f; 14'h2699: x = 16'h202e; 14'h269a: x = 16'h202d; 14'h269b: x = 16'h202c; 14'h269c: x = 16'h202c; 14'h269d: x = 16'h202b; 14'h269e: x = 16'h202a; 14'h269f: x = 16'h2029; 14'h26a0: x = 16'h2028; 14'h26a1: x = 16'h2027; 14'h26a2: x = 16'h2027; 14'h26a3: x = 16'h2026; 14'h26a4: x = 16'h2025; 14'h26a5: x = 16'h2024; 14'h26a6: x = 16'h2023; 14'h26a7: x = 16'h2022; 14'h26a8: x = 16'h2022; 14'h26a9: x = 16'h2021; 14'h26aa: x = 16'h2020; 14'h26ab: x = 16'h201f; 14'h26ac: x = 16'h201e; 14'h26ad: x = 16'h201e; 14'h26ae: x = 16'h201d; 14'h26af: x = 16'h201c; 14'h26b0: x = 16'h201b; 14'h26b1: x = 16'h201a; 14'h26b2: x = 16'h2019; 14'h26b3: x = 16'h2019; 14'h26b4: x = 16'h2018; 14'h26b5: x = 16'h2017; 14'h26b6: x = 16'h2016; 14'h26b7: x = 16'h2015; 14'h26b8: x = 16'h2014; 14'h26b9: x = 16'h2014; 14'h26ba: x = 16'h2013; 14'h26bb: x = 16'h2012; 14'h26bc: x = 16'h2011; 14'h26bd: x = 16'h2010; 14'h26be: x = 16'h200f; 14'h26bf: x = 16'h200f; 14'h26c0: x = 16'h200e; 14'h26c1: x = 16'h200d; 14'h26c2: x = 16'h200c; 14'h26c3: x = 16'h200b; 14'h26c4: x = 16'h200b; 14'h26c5: x = 16'h200a; 14'h26c6: x = 16'h2009; 14'h26c7: x = 16'h2008; 14'h26c8: x = 16'h2007; 14'h26c9: x = 16'h2006; 14'h26ca: x = 16'h2006; 14'h26cb: x = 16'h2005; 14'h26cc: x = 16'h2004; 14'h26cd: x = 16'h2003; 14'h26ce: x = 16'h2002; 14'h26cf: x = 16'h2001; 14'h26d0: x = 16'h2001; 14'h26d1: x = 16'h2000; 14'h26d2: x = 16'h1fff; 14'h26d3: x = 16'h1ffe; 14'h26d4: x = 16'h1ffd; 14'h26d5: x = 16'h1ffd; 14'h26d6: x = 16'h1ffc; 14'h26d7: x = 16'h1ffb; 14'h26d8: x = 16'h1ffa; 14'h26d9: x = 16'h1ff9; 14'h26da: x = 16'h1ff8; 14'h26db: x = 16'h1ff8; 14'h26dc: x = 16'h1ff7; 14'h26dd: x = 16'h1ff6; 14'h26de: x = 16'h1ff5; 14'h26df: x = 16'h1ff4; 14'h26e0: x = 16'h1ff3; 14'h26e1: x = 16'h1ff3; 14'h26e2: x = 16'h1ff2; 14'h26e3: x = 16'h1ff1; 14'h26e4: x = 16'h1ff0; 14'h26e5: x = 16'h1fef; 14'h26e6: x = 16'h1fef; 14'h26e7: x = 16'h1fee; 14'h26e8: x = 16'h1fed; 14'h26e9: x = 16'h1fec; 14'h26ea: x = 16'h1feb; 14'h26eb: x = 16'h1fea; 14'h26ec: x = 16'h1fea; 14'h26ed: x = 16'h1fe9; 14'h26ee: x = 16'h1fe8; 14'h26ef: x = 16'h1fe7; 14'h26f0: x = 16'h1fe6; 14'h26f1: x = 16'h1fe5; 14'h26f2: x = 16'h1fe5; 14'h26f3: x = 16'h1fe4; 14'h26f4: x = 16'h1fe3; 14'h26f5: x = 16'h1fe2; 14'h26f6: x = 16'h1fe1; 14'h26f7: x = 16'h1fe1; 14'h26f8: x = 16'h1fe0; 14'h26f9: x = 16'h1fdf; 14'h26fa: x = 16'h1fde; 14'h26fb: x = 16'h1fdd; 14'h26fc: x = 16'h1fdc; 14'h26fd: x = 16'h1fdc; 14'h26fe: x = 16'h1fdb; 14'h26ff: x = 16'h1fda; 14'h2700: x = 16'h1fd9; 14'h2701: x = 16'h1fd8; 14'h2702: x = 16'h1fd7; 14'h2703: x = 16'h1fd7; 14'h2704: x = 16'h1fd6; 14'h2705: x = 16'h1fd5; 14'h2706: x = 16'h1fd4; 14'h2707: x = 16'h1fd3; 14'h2708: x = 16'h1fd2; 14'h2709: x = 16'h1fd2; 14'h270a: x = 16'h1fd1; 14'h270b: x = 16'h1fd0; 14'h270c: x = 16'h1fcf; 14'h270d: x = 16'h1fce; 14'h270e: x = 16'h1fce; 14'h270f: x = 16'h1fcd; 14'h2710: x = 16'h1fcc; 14'h2711: x = 16'h1fcb; 14'h2712: x = 16'h1fca; 14'h2713: x = 16'h1fc9; 14'h2714: x = 16'h1fc9; 14'h2715: x = 16'h1fc8; 14'h2716: x = 16'h1fc7; 14'h2717: x = 16'h1fc6; 14'h2718: x = 16'h1fc5; 14'h2719: x = 16'h1fc4; 14'h271a: x = 16'h1fc4; 14'h271b: x = 16'h1fc3; 14'h271c: x = 16'h1fc2; 14'h271d: x = 16'h1fc1; 14'h271e: x = 16'h1fc0; 14'h271f: x = 16'h1fc0; 14'h2720: x = 16'h1fbf; 14'h2721: x = 16'h1fbe; 14'h2722: x = 16'h1fbd; 14'h2723: x = 16'h1fbc; 14'h2724: x = 16'h1fbb; 14'h2725: x = 16'h1fbb; 14'h2726: x = 16'h1fba; 14'h2727: x = 16'h1fb9; 14'h2728: x = 16'h1fb8; 14'h2729: x = 16'h1fb7; 14'h272a: x = 16'h1fb6; 14'h272b: x = 16'h1fb6; 14'h272c: x = 16'h1fb5; 14'h272d: x = 16'h1fb4; 14'h272e: x = 16'h1fb3; 14'h272f: x = 16'h1fb2; 14'h2730: x = 16'h1fb2; 14'h2731: x = 16'h1fb1; 14'h2732: x = 16'h1fb0; 14'h2733: x = 16'h1faf; 14'h2734: x = 16'h1fae; 14'h2735: x = 16'h1fad; 14'h2736: x = 16'h1fad; 14'h2737: x = 16'h1fac; 14'h2738: x = 16'h1fab; 14'h2739: x = 16'h1faa; 14'h273a: x = 16'h1fa9; 14'h273b: x = 16'h1fa8; 14'h273c: x = 16'h1fa8; 14'h273d: x = 16'h1fa7; 14'h273e: x = 16'h1fa6; 14'h273f: x = 16'h1fa5; 14'h2740: x = 16'h1fa4; 14'h2741: x = 16'h1fa3; 14'h2742: x = 16'h1fa3; 14'h2743: x = 16'h1fa2; 14'h2744: x = 16'h1fa1; 14'h2745: x = 16'h1fa0; 14'h2746: x = 16'h1f9f; 14'h2747: x = 16'h1f9f; 14'h2748: x = 16'h1f9e; 14'h2749: x = 16'h1f9d; 14'h274a: x = 16'h1f9c; 14'h274b: x = 16'h1f9b; 14'h274c: x = 16'h1f9a; 14'h274d: x = 16'h1f9a; 14'h274e: x = 16'h1f99; 14'h274f: x = 16'h1f98; 14'h2750: x = 16'h1f97; 14'h2751: x = 16'h1f96; 14'h2752: x = 16'h1f95; 14'h2753: x = 16'h1f95; 14'h2754: x = 16'h1f94; 14'h2755: x = 16'h1f93; 14'h2756: x = 16'h1f92; 14'h2757: x = 16'h1f91; 14'h2758: x = 16'h1f91; 14'h2759: x = 16'h1f90; 14'h275a: x = 16'h1f8f; 14'h275b: x = 16'h1f8e; 14'h275c: x = 16'h1f8d; 14'h275d: x = 16'h1f8c; 14'h275e: x = 16'h1f8c; 14'h275f: x = 16'h1f8b; 14'h2760: x = 16'h1f8a; 14'h2761: x = 16'h1f89; 14'h2762: x = 16'h1f88; 14'h2763: x = 16'h1f87; 14'h2764: x = 16'h1f87; 14'h2765: x = 16'h1f86; 14'h2766: x = 16'h1f85; 14'h2767: x = 16'h1f84; 14'h2768: x = 16'h1f83; 14'h2769: x = 16'h1f83; 14'h276a: x = 16'h1f82; 14'h276b: x = 16'h1f81; 14'h276c: x = 16'h1f80; 14'h276d: x = 16'h1f7f; 14'h276e: x = 16'h1f7e; 14'h276f: x = 16'h1f7e; 14'h2770: x = 16'h1f7d; 14'h2771: x = 16'h1f7c; 14'h2772: x = 16'h1f7b; 14'h2773: x = 16'h1f7a; 14'h2774: x = 16'h1f79; 14'h2775: x = 16'h1f79; 14'h2776: x = 16'h1f78; 14'h2777: x = 16'h1f77; 14'h2778: x = 16'h1f76; 14'h2779: x = 16'h1f75; 14'h277a: x = 16'h1f74; 14'h277b: x = 16'h1f74; 14'h277c: x = 16'h1f73; 14'h277d: x = 16'h1f72; 14'h277e: x = 16'h1f71; 14'h277f: x = 16'h1f70; 14'h2780: x = 16'h1f70; 14'h2781: x = 16'h1f6f; 14'h2782: x = 16'h1f6e; 14'h2783: x = 16'h1f6d; 14'h2784: x = 16'h1f6c; 14'h2785: x = 16'h1f6b; 14'h2786: x = 16'h1f6b; 14'h2787: x = 16'h1f6a; 14'h2788: x = 16'h1f69; 14'h2789: x = 16'h1f68; 14'h278a: x = 16'h1f67; 14'h278b: x = 16'h1f66; 14'h278c: x = 16'h1f66; 14'h278d: x = 16'h1f65; 14'h278e: x = 16'h1f64; 14'h278f: x = 16'h1f63; 14'h2790: x = 16'h1f62; 14'h2791: x = 16'h1f62; 14'h2792: x = 16'h1f61; 14'h2793: x = 16'h1f60; 14'h2794: x = 16'h1f5f; 14'h2795: x = 16'h1f5e; 14'h2796: x = 16'h1f5d; 14'h2797: x = 16'h1f5d; 14'h2798: x = 16'h1f5c; 14'h2799: x = 16'h1f5b; 14'h279a: x = 16'h1f5a; 14'h279b: x = 16'h1f59; 14'h279c: x = 16'h1f58; 14'h279d: x = 16'h1f58; 14'h279e: x = 16'h1f57; 14'h279f: x = 16'h1f56; 14'h27a0: x = 16'h1f55; 14'h27a1: x = 16'h1f54; 14'h27a2: x = 16'h1f54; 14'h27a3: x = 16'h1f53; 14'h27a4: x = 16'h1f52; 14'h27a5: x = 16'h1f51; 14'h27a6: x = 16'h1f50; 14'h27a7: x = 16'h1f4f; 14'h27a8: x = 16'h1f4f; 14'h27a9: x = 16'h1f4e; 14'h27aa: x = 16'h1f4d; 14'h27ab: x = 16'h1f4c; 14'h27ac: x = 16'h1f4b; 14'h27ad: x = 16'h1f4a; 14'h27ae: x = 16'h1f4a; 14'h27af: x = 16'h1f49; 14'h27b0: x = 16'h1f48; 14'h27b1: x = 16'h1f47; 14'h27b2: x = 16'h1f46; 14'h27b3: x = 16'h1f45; 14'h27b4: x = 16'h1f45; 14'h27b5: x = 16'h1f44; 14'h27b6: x = 16'h1f43; 14'h27b7: x = 16'h1f42; 14'h27b8: x = 16'h1f41; 14'h27b9: x = 16'h1f41; 14'h27ba: x = 16'h1f40; 14'h27bb: x = 16'h1f3f; 14'h27bc: x = 16'h1f3e; 14'h27bd: x = 16'h1f3d; 14'h27be: x = 16'h1f3c; 14'h27bf: x = 16'h1f3c; 14'h27c0: x = 16'h1f3b; 14'h27c1: x = 16'h1f3a; 14'h27c2: x = 16'h1f39; 14'h27c3: x = 16'h1f38; 14'h27c4: x = 16'h1f37; 14'h27c5: x = 16'h1f37; 14'h27c6: x = 16'h1f36; 14'h27c7: x = 16'h1f35; 14'h27c8: x = 16'h1f34; 14'h27c9: x = 16'h1f33; 14'h27ca: x = 16'h1f33; 14'h27cb: x = 16'h1f32; 14'h27cc: x = 16'h1f31; 14'h27cd: x = 16'h1f30; 14'h27ce: x = 16'h1f2f; 14'h27cf: x = 16'h1f2e; 14'h27d0: x = 16'h1f2e; 14'h27d1: x = 16'h1f2d; 14'h27d2: x = 16'h1f2c; 14'h27d3: x = 16'h1f2b; 14'h27d4: x = 16'h1f2a; 14'h27d5: x = 16'h1f29; 14'h27d6: x = 16'h1f29; 14'h27d7: x = 16'h1f28; 14'h27d8: x = 16'h1f27; 14'h27d9: x = 16'h1f26; 14'h27da: x = 16'h1f25; 14'h27db: x = 16'h1f24; 14'h27dc: x = 16'h1f24; 14'h27dd: x = 16'h1f23; 14'h27de: x = 16'h1f22; 14'h27df: x = 16'h1f21; 14'h27e0: x = 16'h1f20; 14'h27e1: x = 16'h1f20; 14'h27e2: x = 16'h1f1f; 14'h27e3: x = 16'h1f1e; 14'h27e4: x = 16'h1f1d; 14'h27e5: x = 16'h1f1c; 14'h27e6: x = 16'h1f1b; 14'h27e7: x = 16'h1f1b; 14'h27e8: x = 16'h1f1a; 14'h27e9: x = 16'h1f19; 14'h27ea: x = 16'h1f18; 14'h27eb: x = 16'h1f17; 14'h27ec: x = 16'h1f16; 14'h27ed: x = 16'h1f16; 14'h27ee: x = 16'h1f15; 14'h27ef: x = 16'h1f14; 14'h27f0: x = 16'h1f13; 14'h27f1: x = 16'h1f12; 14'h27f2: x = 16'h1f12; 14'h27f3: x = 16'h1f11; 14'h27f4: x = 16'h1f10; 14'h27f5: x = 16'h1f0f; 14'h27f6: x = 16'h1f0e; 14'h27f7: x = 16'h1f0d; 14'h27f8: x = 16'h1f0d; 14'h27f9: x = 16'h1f0c; 14'h27fa: x = 16'h1f0b; 14'h27fb: x = 16'h1f0a; 14'h27fc: x = 16'h1f09; 14'h27fd: x = 16'h1f08; 14'h27fe: x = 16'h1f08; 14'h27ff: x = 16'h1f07; 14'h2800: x = 16'h1f06; 14'h2801: x = 16'h1f05; 14'h2802: x = 16'h1f04; 14'h2803: x = 16'h1f03; 14'h2804: x = 16'h1f03; 14'h2805: x = 16'h1f02; 14'h2806: x = 16'h1f01; 14'h2807: x = 16'h1f00; 14'h2808: x = 16'h1eff; 14'h2809: x = 16'h1eff; 14'h280a: x = 16'h1efe; 14'h280b: x = 16'h1efd; 14'h280c: x = 16'h1efc; 14'h280d: x = 16'h1efb; 14'h280e: x = 16'h1efa; 14'h280f: x = 16'h1efa; 14'h2810: x = 16'h1ef9; 14'h2811: x = 16'h1ef8; 14'h2812: x = 16'h1ef7; 14'h2813: x = 16'h1ef6; 14'h2814: x = 16'h1ef5; 14'h2815: x = 16'h1ef5; 14'h2816: x = 16'h1ef4; 14'h2817: x = 16'h1ef3; 14'h2818: x = 16'h1ef2; 14'h2819: x = 16'h1ef1; 14'h281a: x = 16'h1ef1; 14'h281b: x = 16'h1ef0; 14'h281c: x = 16'h1eef; 14'h281d: x = 16'h1eee; 14'h281e: x = 16'h1eed; 14'h281f: x = 16'h1eec; 14'h2820: x = 16'h1eec; 14'h2821: x = 16'h1eeb; 14'h2822: x = 16'h1eea; 14'h2823: x = 16'h1ee9; 14'h2824: x = 16'h1ee8; 14'h2825: x = 16'h1ee7; 14'h2826: x = 16'h1ee7; 14'h2827: x = 16'h1ee6; 14'h2828: x = 16'h1ee5; 14'h2829: x = 16'h1ee4; 14'h282a: x = 16'h1ee3; 14'h282b: x = 16'h1ee2; 14'h282c: x = 16'h1ee2; 14'h282d: x = 16'h1ee1; 14'h282e: x = 16'h1ee0; 14'h282f: x = 16'h1edf; 14'h2830: x = 16'h1ede; 14'h2831: x = 16'h1ede; 14'h2832: x = 16'h1edd; 14'h2833: x = 16'h1edc; 14'h2834: x = 16'h1edb; 14'h2835: x = 16'h1eda; 14'h2836: x = 16'h1ed9; 14'h2837: x = 16'h1ed9; 14'h2838: x = 16'h1ed8; 14'h2839: x = 16'h1ed7; 14'h283a: x = 16'h1ed6; 14'h283b: x = 16'h1ed5; 14'h283c: x = 16'h1ed4; 14'h283d: x = 16'h1ed4; 14'h283e: x = 16'h1ed3; 14'h283f: x = 16'h1ed2; 14'h2840: x = 16'h1ed1; 14'h2841: x = 16'h1ed0; 14'h2842: x = 16'h1ecf; 14'h2843: x = 16'h1ecf; 14'h2844: x = 16'h1ece; 14'h2845: x = 16'h1ecd; 14'h2846: x = 16'h1ecc; 14'h2847: x = 16'h1ecb; 14'h2848: x = 16'h1ecb; 14'h2849: x = 16'h1eca; 14'h284a: x = 16'h1ec9; 14'h284b: x = 16'h1ec8; 14'h284c: x = 16'h1ec7; 14'h284d: x = 16'h1ec6; 14'h284e: x = 16'h1ec6; 14'h284f: x = 16'h1ec5; 14'h2850: x = 16'h1ec4; 14'h2851: x = 16'h1ec3; 14'h2852: x = 16'h1ec2; 14'h2853: x = 16'h1ec1; 14'h2854: x = 16'h1ec1; 14'h2855: x = 16'h1ec0; 14'h2856: x = 16'h1ebf; 14'h2857: x = 16'h1ebe; 14'h2858: x = 16'h1ebd; 14'h2859: x = 16'h1ebd; 14'h285a: x = 16'h1ebc; 14'h285b: x = 16'h1ebb; 14'h285c: x = 16'h1eba; 14'h285d: x = 16'h1eb9; 14'h285e: x = 16'h1eb8; 14'h285f: x = 16'h1eb8; 14'h2860: x = 16'h1eb7; 14'h2861: x = 16'h1eb6; 14'h2862: x = 16'h1eb5; 14'h2863: x = 16'h1eb4; 14'h2864: x = 16'h1eb3; 14'h2865: x = 16'h1eb3; 14'h2866: x = 16'h1eb2; 14'h2867: x = 16'h1eb1; 14'h2868: x = 16'h1eb0; 14'h2869: x = 16'h1eaf; 14'h286a: x = 16'h1eae; 14'h286b: x = 16'h1eae; 14'h286c: x = 16'h1ead; 14'h286d: x = 16'h1eac; 14'h286e: x = 16'h1eab; 14'h286f: x = 16'h1eaa; 14'h2870: x = 16'h1eaa; 14'h2871: x = 16'h1ea9; 14'h2872: x = 16'h1ea8; 14'h2873: x = 16'h1ea7; 14'h2874: x = 16'h1ea6; 14'h2875: x = 16'h1ea5; 14'h2876: x = 16'h1ea5; 14'h2877: x = 16'h1ea4; 14'h2878: x = 16'h1ea3; 14'h2879: x = 16'h1ea2; 14'h287a: x = 16'h1ea1; 14'h287b: x = 16'h1ea0; 14'h287c: x = 16'h1ea0; 14'h287d: x = 16'h1e9f; 14'h287e: x = 16'h1e9e; 14'h287f: x = 16'h1e9d; 14'h2880: x = 16'h1e9c; 14'h2881: x = 16'h1e9b; 14'h2882: x = 16'h1e9b; 14'h2883: x = 16'h1e9a; 14'h2884: x = 16'h1e99; 14'h2885: x = 16'h1e98; 14'h2886: x = 16'h1e97; 14'h2887: x = 16'h1e97; 14'h2888: x = 16'h1e96; 14'h2889: x = 16'h1e95; 14'h288a: x = 16'h1e94; 14'h288b: x = 16'h1e93; 14'h288c: x = 16'h1e92; 14'h288d: x = 16'h1e92; 14'h288e: x = 16'h1e91; 14'h288f: x = 16'h1e90; 14'h2890: x = 16'h1e8f; 14'h2891: x = 16'h1e8e; 14'h2892: x = 16'h1e8d; 14'h2893: x = 16'h1e8d; 14'h2894: x = 16'h1e8c; 14'h2895: x = 16'h1e8b; 14'h2896: x = 16'h1e8a; 14'h2897: x = 16'h1e89; 14'h2898: x = 16'h1e88; 14'h2899: x = 16'h1e88; 14'h289a: x = 16'h1e87; 14'h289b: x = 16'h1e86; 14'h289c: x = 16'h1e85; 14'h289d: x = 16'h1e84; 14'h289e: x = 16'h1e84; 14'h289f: x = 16'h1e83; 14'h28a0: x = 16'h1e82; 14'h28a1: x = 16'h1e81; 14'h28a2: x = 16'h1e80; 14'h28a3: x = 16'h1e7f; 14'h28a4: x = 16'h1e7f; 14'h28a5: x = 16'h1e7e; 14'h28a6: x = 16'h1e7d; 14'h28a7: x = 16'h1e7c; 14'h28a8: x = 16'h1e7b; 14'h28a9: x = 16'h1e7a; 14'h28aa: x = 16'h1e7a; 14'h28ab: x = 16'h1e79; 14'h28ac: x = 16'h1e78; 14'h28ad: x = 16'h1e77; 14'h28ae: x = 16'h1e76; 14'h28af: x = 16'h1e75; 14'h28b0: x = 16'h1e75; 14'h28b1: x = 16'h1e74; 14'h28b2: x = 16'h1e73; 14'h28b3: x = 16'h1e72; 14'h28b4: x = 16'h1e71; 14'h28b5: x = 16'h1e71; 14'h28b6: x = 16'h1e70; 14'h28b7: x = 16'h1e6f; 14'h28b8: x = 16'h1e6e; 14'h28b9: x = 16'h1e6d; 14'h28ba: x = 16'h1e6c; 14'h28bb: x = 16'h1e6c; 14'h28bc: x = 16'h1e6b; 14'h28bd: x = 16'h1e6a; 14'h28be: x = 16'h1e69; 14'h28bf: x = 16'h1e68; 14'h28c0: x = 16'h1e67; 14'h28c1: x = 16'h1e67; 14'h28c2: x = 16'h1e66; 14'h28c3: x = 16'h1e65; 14'h28c4: x = 16'h1e64; 14'h28c5: x = 16'h1e63; 14'h28c6: x = 16'h1e62; 14'h28c7: x = 16'h1e62; 14'h28c8: x = 16'h1e61; 14'h28c9: x = 16'h1e60; 14'h28ca: x = 16'h1e5f; 14'h28cb: x = 16'h1e5e; 14'h28cc: x = 16'h1e5e; 14'h28cd: x = 16'h1e5d; 14'h28ce: x = 16'h1e5c; 14'h28cf: x = 16'h1e5b; 14'h28d0: x = 16'h1e5a; 14'h28d1: x = 16'h1e59; 14'h28d2: x = 16'h1e59; 14'h28d3: x = 16'h1e58; 14'h28d4: x = 16'h1e57; 14'h28d5: x = 16'h1e56; 14'h28d6: x = 16'h1e55; 14'h28d7: x = 16'h1e54; 14'h28d8: x = 16'h1e54; 14'h28d9: x = 16'h1e53; 14'h28da: x = 16'h1e52; 14'h28db: x = 16'h1e51; 14'h28dc: x = 16'h1e50; 14'h28dd: x = 16'h1e4f; 14'h28de: x = 16'h1e4f; 14'h28df: x = 16'h1e4e; 14'h28e0: x = 16'h1e4d; 14'h28e1: x = 16'h1e4c; 14'h28e2: x = 16'h1e4b; 14'h28e3: x = 16'h1e4a; 14'h28e4: x = 16'h1e4a; 14'h28e5: x = 16'h1e49; 14'h28e6: x = 16'h1e48; 14'h28e7: x = 16'h1e47; 14'h28e8: x = 16'h1e46; 14'h28e9: x = 16'h1e46; 14'h28ea: x = 16'h1e45; 14'h28eb: x = 16'h1e44; 14'h28ec: x = 16'h1e43; 14'h28ed: x = 16'h1e42; 14'h28ee: x = 16'h1e41; 14'h28ef: x = 16'h1e41; 14'h28f0: x = 16'h1e40; 14'h28f1: x = 16'h1e3f; 14'h28f2: x = 16'h1e3e; 14'h28f3: x = 16'h1e3d; 14'h28f4: x = 16'h1e3c; 14'h28f5: x = 16'h1e3c; 14'h28f6: x = 16'h1e3b; 14'h28f7: x = 16'h1e3a; 14'h28f8: x = 16'h1e39; 14'h28f9: x = 16'h1e38; 14'h28fa: x = 16'h1e37; 14'h28fb: x = 16'h1e37; 14'h28fc: x = 16'h1e36; 14'h28fd: x = 16'h1e35; 14'h28fe: x = 16'h1e34; 14'h28ff: x = 16'h1e33; 14'h2900: x = 16'h1e33; 14'h2901: x = 16'h1e32; 14'h2902: x = 16'h1e31; 14'h2903: x = 16'h1e30; 14'h2904: x = 16'h1e2f; 14'h2905: x = 16'h1e2e; 14'h2906: x = 16'h1e2e; 14'h2907: x = 16'h1e2d; 14'h2908: x = 16'h1e2c; 14'h2909: x = 16'h1e2b; 14'h290a: x = 16'h1e2a; 14'h290b: x = 16'h1e29; 14'h290c: x = 16'h1e29; 14'h290d: x = 16'h1e28; 14'h290e: x = 16'h1e27; 14'h290f: x = 16'h1e26; 14'h2910: x = 16'h1e25; 14'h2911: x = 16'h1e24; 14'h2912: x = 16'h1e24; 14'h2913: x = 16'h1e23; 14'h2914: x = 16'h1e22; 14'h2915: x = 16'h1e21; 14'h2916: x = 16'h1e20; 14'h2917: x = 16'h1e1f; 14'h2918: x = 16'h1e1f; 14'h2919: x = 16'h1e1e; 14'h291a: x = 16'h1e1d; 14'h291b: x = 16'h1e1c; 14'h291c: x = 16'h1e1b; 14'h291d: x = 16'h1e1b; 14'h291e: x = 16'h1e1a; 14'h291f: x = 16'h1e19; 14'h2920: x = 16'h1e18; 14'h2921: x = 16'h1e17; 14'h2922: x = 16'h1e16; 14'h2923: x = 16'h1e16; 14'h2924: x = 16'h1e15; 14'h2925: x = 16'h1e14; 14'h2926: x = 16'h1e13; 14'h2927: x = 16'h1e12; 14'h2928: x = 16'h1e11; 14'h2929: x = 16'h1e11; 14'h292a: x = 16'h1e10; 14'h292b: x = 16'h1e0f; 14'h292c: x = 16'h1e0e; 14'h292d: x = 16'h1e0d; 14'h292e: x = 16'h1e0c; 14'h292f: x = 16'h1e0c; 14'h2930: x = 16'h1e0b; 14'h2931: x = 16'h1e0a; 14'h2932: x = 16'h1e09; 14'h2933: x = 16'h1e08; 14'h2934: x = 16'h1e07; 14'h2935: x = 16'h1e07; 14'h2936: x = 16'h1e06; 14'h2937: x = 16'h1e05; 14'h2938: x = 16'h1e04; 14'h2939: x = 16'h1e03; 14'h293a: x = 16'h1e03; 14'h293b: x = 16'h1e02; 14'h293c: x = 16'h1e01; 14'h293d: x = 16'h1e00; 14'h293e: x = 16'h1dff; 14'h293f: x = 16'h1dfe; 14'h2940: x = 16'h1dfe; 14'h2941: x = 16'h1dfd; 14'h2942: x = 16'h1dfc; 14'h2943: x = 16'h1dfb; 14'h2944: x = 16'h1dfa; 14'h2945: x = 16'h1df9; 14'h2946: x = 16'h1df9; 14'h2947: x = 16'h1df8; 14'h2948: x = 16'h1df7; 14'h2949: x = 16'h1df6; 14'h294a: x = 16'h1df5; 14'h294b: x = 16'h1df4; 14'h294c: x = 16'h1df4; 14'h294d: x = 16'h1df3; 14'h294e: x = 16'h1df2; 14'h294f: x = 16'h1df1; 14'h2950: x = 16'h1df0; 14'h2951: x = 16'h1def; 14'h2952: x = 16'h1def; 14'h2953: x = 16'h1dee; 14'h2954: x = 16'h1ded; 14'h2955: x = 16'h1dec; 14'h2956: x = 16'h1deb; 14'h2957: x = 16'h1deb; 14'h2958: x = 16'h1dea; 14'h2959: x = 16'h1de9; 14'h295a: x = 16'h1de8; 14'h295b: x = 16'h1de7; 14'h295c: x = 16'h1de6; 14'h295d: x = 16'h1de6; 14'h295e: x = 16'h1de5; 14'h295f: x = 16'h1de4; 14'h2960: x = 16'h1de3; 14'h2961: x = 16'h1de2; 14'h2962: x = 16'h1de1; 14'h2963: x = 16'h1de1; 14'h2964: x = 16'h1de0; 14'h2965: x = 16'h1ddf; 14'h2966: x = 16'h1dde; 14'h2967: x = 16'h1ddd; 14'h2968: x = 16'h1ddc; 14'h2969: x = 16'h1ddc; 14'h296a: x = 16'h1ddb; 14'h296b: x = 16'h1dda; 14'h296c: x = 16'h1dd9; 14'h296d: x = 16'h1dd8; 14'h296e: x = 16'h1dd7; 14'h296f: x = 16'h1dd7; 14'h2970: x = 16'h1dd6; 14'h2971: x = 16'h1dd5; 14'h2972: x = 16'h1dd4; 14'h2973: x = 16'h1dd3; 14'h2974: x = 16'h1dd3; 14'h2975: x = 16'h1dd2; 14'h2976: x = 16'h1dd1; 14'h2977: x = 16'h1dd0; 14'h2978: x = 16'h1dcf; 14'h2979: x = 16'h1dce; 14'h297a: x = 16'h1dce; 14'h297b: x = 16'h1dcd; 14'h297c: x = 16'h1dcc; 14'h297d: x = 16'h1dcb; 14'h297e: x = 16'h1dca; 14'h297f: x = 16'h1dc9; 14'h2980: x = 16'h1dc9; 14'h2981: x = 16'h1dc8; 14'h2982: x = 16'h1dc7; 14'h2983: x = 16'h1dc6; 14'h2984: x = 16'h1dc5; 14'h2985: x = 16'h1dc4; 14'h2986: x = 16'h1dc4; 14'h2987: x = 16'h1dc3; 14'h2988: x = 16'h1dc2; 14'h2989: x = 16'h1dc1; 14'h298a: x = 16'h1dc0; 14'h298b: x = 16'h1dbf; 14'h298c: x = 16'h1dbf; 14'h298d: x = 16'h1dbe; 14'h298e: x = 16'h1dbd; 14'h298f: x = 16'h1dbc; 14'h2990: x = 16'h1dbb; 14'h2991: x = 16'h1dba; 14'h2992: x = 16'h1dba; 14'h2993: x = 16'h1db9; 14'h2994: x = 16'h1db8; 14'h2995: x = 16'h1db7; 14'h2996: x = 16'h1db6; 14'h2997: x = 16'h1db6; 14'h2998: x = 16'h1db5; 14'h2999: x = 16'h1db4; 14'h299a: x = 16'h1db3; 14'h299b: x = 16'h1db2; 14'h299c: x = 16'h1db1; 14'h299d: x = 16'h1db1; 14'h299e: x = 16'h1db0; 14'h299f: x = 16'h1daf; 14'h29a0: x = 16'h1dae; 14'h29a1: x = 16'h1dad; 14'h29a2: x = 16'h1dac; 14'h29a3: x = 16'h1dac; 14'h29a4: x = 16'h1dab; 14'h29a5: x = 16'h1daa; 14'h29a6: x = 16'h1da9; 14'h29a7: x = 16'h1da8; 14'h29a8: x = 16'h1da7; 14'h29a9: x = 16'h1da7; 14'h29aa: x = 16'h1da6; 14'h29ab: x = 16'h1da5; 14'h29ac: x = 16'h1da4; 14'h29ad: x = 16'h1da3; 14'h29ae: x = 16'h1da2; 14'h29af: x = 16'h1da2; 14'h29b0: x = 16'h1da1; 14'h29b1: x = 16'h1da0; 14'h29b2: x = 16'h1d9f; 14'h29b3: x = 16'h1d9e; 14'h29b4: x = 16'h1d9d; 14'h29b5: x = 16'h1d9d; 14'h29b6: x = 16'h1d9c; 14'h29b7: x = 16'h1d9b; 14'h29b8: x = 16'h1d9a; 14'h29b9: x = 16'h1d99; 14'h29ba: x = 16'h1d99; 14'h29bb: x = 16'h1d98; 14'h29bc: x = 16'h1d97; 14'h29bd: x = 16'h1d96; 14'h29be: x = 16'h1d95; 14'h29bf: x = 16'h1d94; 14'h29c0: x = 16'h1d94; 14'h29c1: x = 16'h1d93; 14'h29c2: x = 16'h1d92; 14'h29c3: x = 16'h1d91; 14'h29c4: x = 16'h1d90; 14'h29c5: x = 16'h1d8f; 14'h29c6: x = 16'h1d8f; 14'h29c7: x = 16'h1d8e; 14'h29c8: x = 16'h1d8d; 14'h29c9: x = 16'h1d8c; 14'h29ca: x = 16'h1d8b; 14'h29cb: x = 16'h1d8a; 14'h29cc: x = 16'h1d8a; 14'h29cd: x = 16'h1d89; 14'h29ce: x = 16'h1d88; 14'h29cf: x = 16'h1d87; 14'h29d0: x = 16'h1d86; 14'h29d1: x = 16'h1d85; 14'h29d2: x = 16'h1d85; 14'h29d3: x = 16'h1d84; 14'h29d4: x = 16'h1d83; 14'h29d5: x = 16'h1d82; 14'h29d6: x = 16'h1d81; 14'h29d7: x = 16'h1d80; 14'h29d8: x = 16'h1d80; 14'h29d9: x = 16'h1d7f; 14'h29da: x = 16'h1d7e; 14'h29db: x = 16'h1d7d; 14'h29dc: x = 16'h1d7c; 14'h29dd: x = 16'h1d7b; 14'h29de: x = 16'h1d7b; 14'h29df: x = 16'h1d7a; 14'h29e0: x = 16'h1d79; 14'h29e1: x = 16'h1d78; 14'h29e2: x = 16'h1d77; 14'h29e3: x = 16'h1d76; 14'h29e4: x = 16'h1d76; 14'h29e5: x = 16'h1d75; 14'h29e6: x = 16'h1d74; 14'h29e7: x = 16'h1d73; 14'h29e8: x = 16'h1d72; 14'h29e9: x = 16'h1d72; 14'h29ea: x = 16'h1d71; 14'h29eb: x = 16'h1d70; 14'h29ec: x = 16'h1d6f; 14'h29ed: x = 16'h1d6e; 14'h29ee: x = 16'h1d6d; 14'h29ef: x = 16'h1d6d; 14'h29f0: x = 16'h1d6c; 14'h29f1: x = 16'h1d6b; 14'h29f2: x = 16'h1d6a; 14'h29f3: x = 16'h1d69; 14'h29f4: x = 16'h1d68; 14'h29f5: x = 16'h1d68; 14'h29f6: x = 16'h1d67; 14'h29f7: x = 16'h1d66; 14'h29f8: x = 16'h1d65; 14'h29f9: x = 16'h1d64; 14'h29fa: x = 16'h1d63; 14'h29fb: x = 16'h1d63; 14'h29fc: x = 16'h1d62; 14'h29fd: x = 16'h1d61; 14'h29fe: x = 16'h1d60; 14'h29ff: x = 16'h1d5f; 14'h2a00: x = 16'h1d5e; 14'h2a01: x = 16'h1d5e; 14'h2a02: x = 16'h1d5d; 14'h2a03: x = 16'h1d5c; 14'h2a04: x = 16'h1d5b; 14'h2a05: x = 16'h1d5a; 14'h2a06: x = 16'h1d59; 14'h2a07: x = 16'h1d59; 14'h2a08: x = 16'h1d58; 14'h2a09: x = 16'h1d57; 14'h2a0a: x = 16'h1d56; 14'h2a0b: x = 16'h1d55; 14'h2a0c: x = 16'h1d54; 14'h2a0d: x = 16'h1d54; 14'h2a0e: x = 16'h1d53; 14'h2a0f: x = 16'h1d52; 14'h2a10: x = 16'h1d51; 14'h2a11: x = 16'h1d50; 14'h2a12: x = 16'h1d4f; 14'h2a13: x = 16'h1d4f; 14'h2a14: x = 16'h1d4e; 14'h2a15: x = 16'h1d4d; 14'h2a16: x = 16'h1d4c; 14'h2a17: x = 16'h1d4b; 14'h2a18: x = 16'h1d4b; 14'h2a19: x = 16'h1d4a; 14'h2a1a: x = 16'h1d49; 14'h2a1b: x = 16'h1d48; 14'h2a1c: x = 16'h1d47; 14'h2a1d: x = 16'h1d46; 14'h2a1e: x = 16'h1d46; 14'h2a1f: x = 16'h1d45; 14'h2a20: x = 16'h1d44; 14'h2a21: x = 16'h1d43; 14'h2a22: x = 16'h1d42; 14'h2a23: x = 16'h1d41; 14'h2a24: x = 16'h1d41; 14'h2a25: x = 16'h1d40; 14'h2a26: x = 16'h1d3f; 14'h2a27: x = 16'h1d3e; 14'h2a28: x = 16'h1d3d; 14'h2a29: x = 16'h1d3c; 14'h2a2a: x = 16'h1d3c; 14'h2a2b: x = 16'h1d3b; 14'h2a2c: x = 16'h1d3a; 14'h2a2d: x = 16'h1d39; 14'h2a2e: x = 16'h1d38; 14'h2a2f: x = 16'h1d37; 14'h2a30: x = 16'h1d37; 14'h2a31: x = 16'h1d36; 14'h2a32: x = 16'h1d35; 14'h2a33: x = 16'h1d34; 14'h2a34: x = 16'h1d33; 14'h2a35: x = 16'h1d32; 14'h2a36: x = 16'h1d32; 14'h2a37: x = 16'h1d31; 14'h2a38: x = 16'h1d30; 14'h2a39: x = 16'h1d2f; 14'h2a3a: x = 16'h1d2e; 14'h2a3b: x = 16'h1d2d; 14'h2a3c: x = 16'h1d2d; 14'h2a3d: x = 16'h1d2c; 14'h2a3e: x = 16'h1d2b; 14'h2a3f: x = 16'h1d2a; 14'h2a40: x = 16'h1d29; 14'h2a41: x = 16'h1d28; 14'h2a42: x = 16'h1d28; 14'h2a43: x = 16'h1d27; 14'h2a44: x = 16'h1d26; 14'h2a45: x = 16'h1d25; 14'h2a46: x = 16'h1d24; 14'h2a47: x = 16'h1d23; 14'h2a48: x = 16'h1d23; 14'h2a49: x = 16'h1d22; 14'h2a4a: x = 16'h1d21; 14'h2a4b: x = 16'h1d20; 14'h2a4c: x = 16'h1d1f; 14'h2a4d: x = 16'h1d1e; 14'h2a4e: x = 16'h1d1e; 14'h2a4f: x = 16'h1d1d; 14'h2a50: x = 16'h1d1c; 14'h2a51: x = 16'h1d1b; 14'h2a52: x = 16'h1d1a; 14'h2a53: x = 16'h1d19; 14'h2a54: x = 16'h1d19; 14'h2a55: x = 16'h1d18; 14'h2a56: x = 16'h1d17; 14'h2a57: x = 16'h1d16; 14'h2a58: x = 16'h1d15; 14'h2a59: x = 16'h1d14; 14'h2a5a: x = 16'h1d14; 14'h2a5b: x = 16'h1d13; 14'h2a5c: x = 16'h1d12; 14'h2a5d: x = 16'h1d11; 14'h2a5e: x = 16'h1d10; 14'h2a5f: x = 16'h1d10; 14'h2a60: x = 16'h1d0f; 14'h2a61: x = 16'h1d0e; 14'h2a62: x = 16'h1d0d; 14'h2a63: x = 16'h1d0c; 14'h2a64: x = 16'h1d0b; 14'h2a65: x = 16'h1d0b; 14'h2a66: x = 16'h1d0a; 14'h2a67: x = 16'h1d09; 14'h2a68: x = 16'h1d08; 14'h2a69: x = 16'h1d07; 14'h2a6a: x = 16'h1d06; 14'h2a6b: x = 16'h1d06; 14'h2a6c: x = 16'h1d05; 14'h2a6d: x = 16'h1d04; 14'h2a6e: x = 16'h1d03; 14'h2a6f: x = 16'h1d02; 14'h2a70: x = 16'h1d01; 14'h2a71: x = 16'h1d01; 14'h2a72: x = 16'h1d00; 14'h2a73: x = 16'h1cff; 14'h2a74: x = 16'h1cfe; 14'h2a75: x = 16'h1cfd; 14'h2a76: x = 16'h1cfc; 14'h2a77: x = 16'h1cfc; 14'h2a78: x = 16'h1cfb; 14'h2a79: x = 16'h1cfa; 14'h2a7a: x = 16'h1cf9; 14'h2a7b: x = 16'h1cf8; 14'h2a7c: x = 16'h1cf7; 14'h2a7d: x = 16'h1cf7; 14'h2a7e: x = 16'h1cf6; 14'h2a7f: x = 16'h1cf5; 14'h2a80: x = 16'h1cf4; 14'h2a81: x = 16'h1cf3; 14'h2a82: x = 16'h1cf2; 14'h2a83: x = 16'h1cf2; 14'h2a84: x = 16'h1cf1; 14'h2a85: x = 16'h1cf0; 14'h2a86: x = 16'h1cef; 14'h2a87: x = 16'h1cee; 14'h2a88: x = 16'h1ced; 14'h2a89: x = 16'h1ced; 14'h2a8a: x = 16'h1cec; 14'h2a8b: x = 16'h1ceb; 14'h2a8c: x = 16'h1cea; 14'h2a8d: x = 16'h1ce9; 14'h2a8e: x = 16'h1ce8; 14'h2a8f: x = 16'h1ce8; 14'h2a90: x = 16'h1ce7; 14'h2a91: x = 16'h1ce6; 14'h2a92: x = 16'h1ce5; 14'h2a93: x = 16'h1ce4; 14'h2a94: x = 16'h1ce3; 14'h2a95: x = 16'h1ce3; 14'h2a96: x = 16'h1ce2; 14'h2a97: x = 16'h1ce1; 14'h2a98: x = 16'h1ce0; 14'h2a99: x = 16'h1cdf; 14'h2a9a: x = 16'h1cde; 14'h2a9b: x = 16'h1cde; 14'h2a9c: x = 16'h1cdd; 14'h2a9d: x = 16'h1cdc; 14'h2a9e: x = 16'h1cdb; 14'h2a9f: x = 16'h1cda; 14'h2aa0: x = 16'h1cd9; 14'h2aa1: x = 16'h1cd9; 14'h2aa2: x = 16'h1cd8; 14'h2aa3: x = 16'h1cd7; 14'h2aa4: x = 16'h1cd6; 14'h2aa5: x = 16'h1cd5; 14'h2aa6: x = 16'h1cd4; 14'h2aa7: x = 16'h1cd4; 14'h2aa8: x = 16'h1cd3; 14'h2aa9: x = 16'h1cd2; 14'h2aaa: x = 16'h1cd1; 14'h2aab: x = 16'h1cd0; 14'h2aac: x = 16'h1ccf; 14'h2aad: x = 16'h1ccf; 14'h2aae: x = 16'h1cce; 14'h2aaf: x = 16'h1ccd; 14'h2ab0: x = 16'h1ccc; 14'h2ab1: x = 16'h1ccb; 14'h2ab2: x = 16'h1cca; 14'h2ab3: x = 16'h1cca; 14'h2ab4: x = 16'h1cc9; 14'h2ab5: x = 16'h1cc8; 14'h2ab6: x = 16'h1cc7; 14'h2ab7: x = 16'h1cc6; 14'h2ab8: x = 16'h1cc5; 14'h2ab9: x = 16'h1cc5; 14'h2aba: x = 16'h1cc4; 14'h2abb: x = 16'h1cc3; 14'h2abc: x = 16'h1cc2; 14'h2abd: x = 16'h1cc1; 14'h2abe: x = 16'h1cc0; 14'h2abf: x = 16'h1cc0; 14'h2ac0: x = 16'h1cbf; 14'h2ac1: x = 16'h1cbe; 14'h2ac2: x = 16'h1cbd; 14'h2ac3: x = 16'h1cbc; 14'h2ac4: x = 16'h1cbb; 14'h2ac5: x = 16'h1cbb; 14'h2ac6: x = 16'h1cba; 14'h2ac7: x = 16'h1cb9; 14'h2ac8: x = 16'h1cb8; 14'h2ac9: x = 16'h1cb7; 14'h2aca: x = 16'h1cb6; 14'h2acb: x = 16'h1cb6; 14'h2acc: x = 16'h1cb5; 14'h2acd: x = 16'h1cb4; 14'h2ace: x = 16'h1cb3; 14'h2acf: x = 16'h1cb2; 14'h2ad0: x = 16'h1cb1; 14'h2ad1: x = 16'h1cb1; 14'h2ad2: x = 16'h1cb0; 14'h2ad3: x = 16'h1caf; 14'h2ad4: x = 16'h1cae; 14'h2ad5: x = 16'h1cad; 14'h2ad6: x = 16'h1cac; 14'h2ad7: x = 16'h1cac; 14'h2ad8: x = 16'h1cab; 14'h2ad9: x = 16'h1caa; 14'h2ada: x = 16'h1ca9; 14'h2adb: x = 16'h1ca8; 14'h2adc: x = 16'h1ca7; 14'h2add: x = 16'h1ca7; 14'h2ade: x = 16'h1ca6; 14'h2adf: x = 16'h1ca5; 14'h2ae0: x = 16'h1ca4; 14'h2ae1: x = 16'h1ca3; 14'h2ae2: x = 16'h1ca2; 14'h2ae3: x = 16'h1ca2; 14'h2ae4: x = 16'h1ca1; 14'h2ae5: x = 16'h1ca0; 14'h2ae6: x = 16'h1c9f; 14'h2ae7: x = 16'h1c9e; 14'h2ae8: x = 16'h1c9d; 14'h2ae9: x = 16'h1c9d; 14'h2aea: x = 16'h1c9c; 14'h2aeb: x = 16'h1c9b; 14'h2aec: x = 16'h1c9a; 14'h2aed: x = 16'h1c99; 14'h2aee: x = 16'h1c98; 14'h2aef: x = 16'h1c98; 14'h2af0: x = 16'h1c97; 14'h2af1: x = 16'h1c96; 14'h2af2: x = 16'h1c95; 14'h2af3: x = 16'h1c94; 14'h2af4: x = 16'h1c93; 14'h2af5: x = 16'h1c93; 14'h2af6: x = 16'h1c92; 14'h2af7: x = 16'h1c91; 14'h2af8: x = 16'h1c90; 14'h2af9: x = 16'h1c8f; 14'h2afa: x = 16'h1c8e; 14'h2afb: x = 16'h1c8e; 14'h2afc: x = 16'h1c8d; 14'h2afd: x = 16'h1c8c; 14'h2afe: x = 16'h1c8b; 14'h2aff: x = 16'h1c8a; 14'h2b00: x = 16'h1c89; 14'h2b01: x = 16'h1c89; 14'h2b02: x = 16'h1c88; 14'h2b03: x = 16'h1c87; 14'h2b04: x = 16'h1c86; 14'h2b05: x = 16'h1c85; 14'h2b06: x = 16'h1c84; 14'h2b07: x = 16'h1c84; 14'h2b08: x = 16'h1c83; 14'h2b09: x = 16'h1c82; 14'h2b0a: x = 16'h1c81; 14'h2b0b: x = 16'h1c80; 14'h2b0c: x = 16'h1c7f; 14'h2b0d: x = 16'h1c7f; 14'h2b0e: x = 16'h1c7e; 14'h2b0f: x = 16'h1c7d; 14'h2b10: x = 16'h1c7c; 14'h2b11: x = 16'h1c7b; 14'h2b12: x = 16'h1c7a; 14'h2b13: x = 16'h1c7a; 14'h2b14: x = 16'h1c79; 14'h2b15: x = 16'h1c78; 14'h2b16: x = 16'h1c77; 14'h2b17: x = 16'h1c76; 14'h2b18: x = 16'h1c75; 14'h2b19: x = 16'h1c75; 14'h2b1a: x = 16'h1c74; 14'h2b1b: x = 16'h1c73; 14'h2b1c: x = 16'h1c72; 14'h2b1d: x = 16'h1c71; 14'h2b1e: x = 16'h1c70; 14'h2b1f: x = 16'h1c70; 14'h2b20: x = 16'h1c6f; 14'h2b21: x = 16'h1c6e; 14'h2b22: x = 16'h1c6d; 14'h2b23: x = 16'h1c6c; 14'h2b24: x = 16'h1c6b; 14'h2b25: x = 16'h1c6b; 14'h2b26: x = 16'h1c6a; 14'h2b27: x = 16'h1c69; 14'h2b28: x = 16'h1c68; 14'h2b29: x = 16'h1c67; 14'h2b2a: x = 16'h1c66; 14'h2b2b: x = 16'h1c65; 14'h2b2c: x = 16'h1c65; 14'h2b2d: x = 16'h1c64; 14'h2b2e: x = 16'h1c63; 14'h2b2f: x = 16'h1c62; 14'h2b30: x = 16'h1c61; 14'h2b31: x = 16'h1c60; 14'h2b32: x = 16'h1c60; 14'h2b33: x = 16'h1c5f; 14'h2b34: x = 16'h1c5e; 14'h2b35: x = 16'h1c5d; 14'h2b36: x = 16'h1c5c; 14'h2b37: x = 16'h1c5b; 14'h2b38: x = 16'h1c5b; 14'h2b39: x = 16'h1c5a; 14'h2b3a: x = 16'h1c59; 14'h2b3b: x = 16'h1c58; 14'h2b3c: x = 16'h1c57; 14'h2b3d: x = 16'h1c56; 14'h2b3e: x = 16'h1c56; 14'h2b3f: x = 16'h1c55; 14'h2b40: x = 16'h1c54; 14'h2b41: x = 16'h1c53; 14'h2b42: x = 16'h1c52; 14'h2b43: x = 16'h1c51; 14'h2b44: x = 16'h1c51; 14'h2b45: x = 16'h1c50; 14'h2b46: x = 16'h1c4f; 14'h2b47: x = 16'h1c4e; 14'h2b48: x = 16'h1c4d; 14'h2b49: x = 16'h1c4c; 14'h2b4a: x = 16'h1c4c; 14'h2b4b: x = 16'h1c4b; 14'h2b4c: x = 16'h1c4a; 14'h2b4d: x = 16'h1c49; 14'h2b4e: x = 16'h1c48; 14'h2b4f: x = 16'h1c47; 14'h2b50: x = 16'h1c47; 14'h2b51: x = 16'h1c46; 14'h2b52: x = 16'h1c45; 14'h2b53: x = 16'h1c44; 14'h2b54: x = 16'h1c43; 14'h2b55: x = 16'h1c42; 14'h2b56: x = 16'h1c42; 14'h2b57: x = 16'h1c41; 14'h2b58: x = 16'h1c40; 14'h2b59: x = 16'h1c3f; 14'h2b5a: x = 16'h1c3e; 14'h2b5b: x = 16'h1c3d; 14'h2b5c: x = 16'h1c3d; 14'h2b5d: x = 16'h1c3c; 14'h2b5e: x = 16'h1c3b; 14'h2b5f: x = 16'h1c3a; 14'h2b60: x = 16'h1c39; 14'h2b61: x = 16'h1c38; 14'h2b62: x = 16'h1c38; 14'h2b63: x = 16'h1c37; 14'h2b64: x = 16'h1c36; 14'h2b65: x = 16'h1c35; 14'h2b66: x = 16'h1c34; 14'h2b67: x = 16'h1c33; 14'h2b68: x = 16'h1c33; 14'h2b69: x = 16'h1c32; 14'h2b6a: x = 16'h1c31; 14'h2b6b: x = 16'h1c30; 14'h2b6c: x = 16'h1c2f; 14'h2b6d: x = 16'h1c2e; 14'h2b6e: x = 16'h1c2d; 14'h2b6f: x = 16'h1c2d; 14'h2b70: x = 16'h1c2c; 14'h2b71: x = 16'h1c2b; 14'h2b72: x = 16'h1c2a; 14'h2b73: x = 16'h1c29; 14'h2b74: x = 16'h1c28; 14'h2b75: x = 16'h1c28; 14'h2b76: x = 16'h1c27; 14'h2b77: x = 16'h1c26; 14'h2b78: x = 16'h1c25; 14'h2b79: x = 16'h1c24; 14'h2b7a: x = 16'h1c23; 14'h2b7b: x = 16'h1c23; 14'h2b7c: x = 16'h1c22; 14'h2b7d: x = 16'h1c21; 14'h2b7e: x = 16'h1c20; 14'h2b7f: x = 16'h1c1f; 14'h2b80: x = 16'h1c1e; 14'h2b81: x = 16'h1c1e; 14'h2b82: x = 16'h1c1d; 14'h2b83: x = 16'h1c1c; 14'h2b84: x = 16'h1c1b; 14'h2b85: x = 16'h1c1a; 14'h2b86: x = 16'h1c19; 14'h2b87: x = 16'h1c19; 14'h2b88: x = 16'h1c18; 14'h2b89: x = 16'h1c17; 14'h2b8a: x = 16'h1c16; 14'h2b8b: x = 16'h1c15; 14'h2b8c: x = 16'h1c14; 14'h2b8d: x = 16'h1c14; 14'h2b8e: x = 16'h1c13; 14'h2b8f: x = 16'h1c12; 14'h2b90: x = 16'h1c11; 14'h2b91: x = 16'h1c10; 14'h2b92: x = 16'h1c0f; 14'h2b93: x = 16'h1c0f; 14'h2b94: x = 16'h1c0e; 14'h2b95: x = 16'h1c0d; 14'h2b96: x = 16'h1c0c; 14'h2b97: x = 16'h1c0b; 14'h2b98: x = 16'h1c0a; 14'h2b99: x = 16'h1c09; 14'h2b9a: x = 16'h1c09; 14'h2b9b: x = 16'h1c08; 14'h2b9c: x = 16'h1c07; 14'h2b9d: x = 16'h1c06; 14'h2b9e: x = 16'h1c05; 14'h2b9f: x = 16'h1c04; 14'h2ba0: x = 16'h1c04; 14'h2ba1: x = 16'h1c03; 14'h2ba2: x = 16'h1c02; 14'h2ba3: x = 16'h1c01; 14'h2ba4: x = 16'h1c00; 14'h2ba5: x = 16'h1bff; 14'h2ba6: x = 16'h1bff; 14'h2ba7: x = 16'h1bfe; 14'h2ba8: x = 16'h1bfd; 14'h2ba9: x = 16'h1bfc; 14'h2baa: x = 16'h1bfb; 14'h2bab: x = 16'h1bfa; 14'h2bac: x = 16'h1bfa; 14'h2bad: x = 16'h1bf9; 14'h2bae: x = 16'h1bf8; 14'h2baf: x = 16'h1bf7; 14'h2bb0: x = 16'h1bf6; 14'h2bb1: x = 16'h1bf5; 14'h2bb2: x = 16'h1bf5; 14'h2bb3: x = 16'h1bf4; 14'h2bb4: x = 16'h1bf3; 14'h2bb5: x = 16'h1bf2; 14'h2bb6: x = 16'h1bf1; 14'h2bb7: x = 16'h1bf0; 14'h2bb8: x = 16'h1bf0; 14'h2bb9: x = 16'h1bef; 14'h2bba: x = 16'h1bee; 14'h2bbb: x = 16'h1bed; 14'h2bbc: x = 16'h1bec; 14'h2bbd: x = 16'h1beb; 14'h2bbe: x = 16'h1bea; 14'h2bbf: x = 16'h1bea; 14'h2bc0: x = 16'h1be9; 14'h2bc1: x = 16'h1be8; 14'h2bc2: x = 16'h1be7; 14'h2bc3: x = 16'h1be6; 14'h2bc4: x = 16'h1be5; 14'h2bc5: x = 16'h1be5; 14'h2bc6: x = 16'h1be4; 14'h2bc7: x = 16'h1be3; 14'h2bc8: x = 16'h1be2; 14'h2bc9: x = 16'h1be1; 14'h2bca: x = 16'h1be0; 14'h2bcb: x = 16'h1be0; 14'h2bcc: x = 16'h1bdf; 14'h2bcd: x = 16'h1bde; 14'h2bce: x = 16'h1bdd; 14'h2bcf: x = 16'h1bdc; 14'h2bd0: x = 16'h1bdb; 14'h2bd1: x = 16'h1bdb; 14'h2bd2: x = 16'h1bda; 14'h2bd3: x = 16'h1bd9; 14'h2bd4: x = 16'h1bd8; 14'h2bd5: x = 16'h1bd7; 14'h2bd6: x = 16'h1bd6; 14'h2bd7: x = 16'h1bd6; 14'h2bd8: x = 16'h1bd5; 14'h2bd9: x = 16'h1bd4; 14'h2bda: x = 16'h1bd3; 14'h2bdb: x = 16'h1bd2; 14'h2bdc: x = 16'h1bd1; 14'h2bdd: x = 16'h1bd0; 14'h2bde: x = 16'h1bd0; 14'h2bdf: x = 16'h1bcf; 14'h2be0: x = 16'h1bce; 14'h2be1: x = 16'h1bcd; 14'h2be2: x = 16'h1bcc; 14'h2be3: x = 16'h1bcb; 14'h2be4: x = 16'h1bcb; 14'h2be5: x = 16'h1bca; 14'h2be6: x = 16'h1bc9; 14'h2be7: x = 16'h1bc8; 14'h2be8: x = 16'h1bc7; 14'h2be9: x = 16'h1bc6; 14'h2bea: x = 16'h1bc6; 14'h2beb: x = 16'h1bc5; 14'h2bec: x = 16'h1bc4; 14'h2bed: x = 16'h1bc3; 14'h2bee: x = 16'h1bc2; 14'h2bef: x = 16'h1bc1; 14'h2bf0: x = 16'h1bc1; 14'h2bf1: x = 16'h1bc0; 14'h2bf2: x = 16'h1bbf; 14'h2bf3: x = 16'h1bbe; 14'h2bf4: x = 16'h1bbd; 14'h2bf5: x = 16'h1bbc; 14'h2bf6: x = 16'h1bbb; 14'h2bf7: x = 16'h1bbb; 14'h2bf8: x = 16'h1bba; 14'h2bf9: x = 16'h1bb9; 14'h2bfa: x = 16'h1bb8; 14'h2bfb: x = 16'h1bb7; 14'h2bfc: x = 16'h1bb6; 14'h2bfd: x = 16'h1bb6; 14'h2bfe: x = 16'h1bb5; 14'h2bff: x = 16'h1bb4; 14'h2c00: x = 16'h1bb3; 14'h2c01: x = 16'h1bb2; 14'h2c02: x = 16'h1bb1; 14'h2c03: x = 16'h1bb1; 14'h2c04: x = 16'h1bb0; 14'h2c05: x = 16'h1baf; 14'h2c06: x = 16'h1bae; 14'h2c07: x = 16'h1bad; 14'h2c08: x = 16'h1bac; 14'h2c09: x = 16'h1bac; 14'h2c0a: x = 16'h1bab; 14'h2c0b: x = 16'h1baa; 14'h2c0c: x = 16'h1ba9; 14'h2c0d: x = 16'h1ba8; 14'h2c0e: x = 16'h1ba7; 14'h2c0f: x = 16'h1ba6; 14'h2c10: x = 16'h1ba6; 14'h2c11: x = 16'h1ba5; 14'h2c12: x = 16'h1ba4; 14'h2c13: x = 16'h1ba3; 14'h2c14: x = 16'h1ba2; 14'h2c15: x = 16'h1ba1; 14'h2c16: x = 16'h1ba1; 14'h2c17: x = 16'h1ba0; 14'h2c18: x = 16'h1b9f; 14'h2c19: x = 16'h1b9e; 14'h2c1a: x = 16'h1b9d; 14'h2c1b: x = 16'h1b9c; 14'h2c1c: x = 16'h1b9c; 14'h2c1d: x = 16'h1b9b; 14'h2c1e: x = 16'h1b9a; 14'h2c1f: x = 16'h1b99; 14'h2c20: x = 16'h1b98; 14'h2c21: x = 16'h1b97; 14'h2c22: x = 16'h1b97; 14'h2c23: x = 16'h1b96; 14'h2c24: x = 16'h1b95; 14'h2c25: x = 16'h1b94; 14'h2c26: x = 16'h1b93; 14'h2c27: x = 16'h1b92; 14'h2c28: x = 16'h1b91; 14'h2c29: x = 16'h1b91; 14'h2c2a: x = 16'h1b90; 14'h2c2b: x = 16'h1b8f; 14'h2c2c: x = 16'h1b8e; 14'h2c2d: x = 16'h1b8d; 14'h2c2e: x = 16'h1b8c; 14'h2c2f: x = 16'h1b8c; 14'h2c30: x = 16'h1b8b; 14'h2c31: x = 16'h1b8a; 14'h2c32: x = 16'h1b89; 14'h2c33: x = 16'h1b88; 14'h2c34: x = 16'h1b87; 14'h2c35: x = 16'h1b87; 14'h2c36: x = 16'h1b86; 14'h2c37: x = 16'h1b85; 14'h2c38: x = 16'h1b84; 14'h2c39: x = 16'h1b83; 14'h2c3a: x = 16'h1b82; 14'h2c3b: x = 16'h1b81; 14'h2c3c: x = 16'h1b81; 14'h2c3d: x = 16'h1b80; 14'h2c3e: x = 16'h1b7f; 14'h2c3f: x = 16'h1b7e; 14'h2c40: x = 16'h1b7d; 14'h2c41: x = 16'h1b7c; 14'h2c42: x = 16'h1b7c; 14'h2c43: x = 16'h1b7b; 14'h2c44: x = 16'h1b7a; 14'h2c45: x = 16'h1b79; 14'h2c46: x = 16'h1b78; 14'h2c47: x = 16'h1b77; 14'h2c48: x = 16'h1b77; 14'h2c49: x = 16'h1b76; 14'h2c4a: x = 16'h1b75; 14'h2c4b: x = 16'h1b74; 14'h2c4c: x = 16'h1b73; 14'h2c4d: x = 16'h1b72; 14'h2c4e: x = 16'h1b71; 14'h2c4f: x = 16'h1b71; 14'h2c50: x = 16'h1b70; 14'h2c51: x = 16'h1b6f; 14'h2c52: x = 16'h1b6e; 14'h2c53: x = 16'h1b6d; 14'h2c54: x = 16'h1b6c; 14'h2c55: x = 16'h1b6c; 14'h2c56: x = 16'h1b6b; 14'h2c57: x = 16'h1b6a; 14'h2c58: x = 16'h1b69; 14'h2c59: x = 16'h1b68; 14'h2c5a: x = 16'h1b67; 14'h2c5b: x = 16'h1b67; 14'h2c5c: x = 16'h1b66; 14'h2c5d: x = 16'h1b65; 14'h2c5e: x = 16'h1b64; 14'h2c5f: x = 16'h1b63; 14'h2c60: x = 16'h1b62; 14'h2c61: x = 16'h1b61; 14'h2c62: x = 16'h1b61; 14'h2c63: x = 16'h1b60; 14'h2c64: x = 16'h1b5f; 14'h2c65: x = 16'h1b5e; 14'h2c66: x = 16'h1b5d; 14'h2c67: x = 16'h1b5c; 14'h2c68: x = 16'h1b5c; 14'h2c69: x = 16'h1b5b; 14'h2c6a: x = 16'h1b5a; 14'h2c6b: x = 16'h1b59; 14'h2c6c: x = 16'h1b58; 14'h2c6d: x = 16'h1b57; 14'h2c6e: x = 16'h1b57; 14'h2c6f: x = 16'h1b56; 14'h2c70: x = 16'h1b55; 14'h2c71: x = 16'h1b54; 14'h2c72: x = 16'h1b53; 14'h2c73: x = 16'h1b52; 14'h2c74: x = 16'h1b51; 14'h2c75: x = 16'h1b51; 14'h2c76: x = 16'h1b50; 14'h2c77: x = 16'h1b4f; 14'h2c78: x = 16'h1b4e; 14'h2c79: x = 16'h1b4d; 14'h2c7a: x = 16'h1b4c; 14'h2c7b: x = 16'h1b4c; 14'h2c7c: x = 16'h1b4b; 14'h2c7d: x = 16'h1b4a; 14'h2c7e: x = 16'h1b49; 14'h2c7f: x = 16'h1b48; 14'h2c80: x = 16'h1b47; 14'h2c81: x = 16'h1b46; 14'h2c82: x = 16'h1b46; 14'h2c83: x = 16'h1b45; 14'h2c84: x = 16'h1b44; 14'h2c85: x = 16'h1b43; 14'h2c86: x = 16'h1b42; 14'h2c87: x = 16'h1b41; 14'h2c88: x = 16'h1b41; 14'h2c89: x = 16'h1b40; 14'h2c8a: x = 16'h1b3f; 14'h2c8b: x = 16'h1b3e; 14'h2c8c: x = 16'h1b3d; 14'h2c8d: x = 16'h1b3c; 14'h2c8e: x = 16'h1b3c; 14'h2c8f: x = 16'h1b3b; 14'h2c90: x = 16'h1b3a; 14'h2c91: x = 16'h1b39; 14'h2c92: x = 16'h1b38; 14'h2c93: x = 16'h1b37; 14'h2c94: x = 16'h1b36; 14'h2c95: x = 16'h1b36; 14'h2c96: x = 16'h1b35; 14'h2c97: x = 16'h1b34; 14'h2c98: x = 16'h1b33; 14'h2c99: x = 16'h1b32; 14'h2c9a: x = 16'h1b31; 14'h2c9b: x = 16'h1b31; 14'h2c9c: x = 16'h1b30; 14'h2c9d: x = 16'h1b2f; 14'h2c9e: x = 16'h1b2e; 14'h2c9f: x = 16'h1b2d; 14'h2ca0: x = 16'h1b2c; 14'h2ca1: x = 16'h1b2b; 14'h2ca2: x = 16'h1b2b; 14'h2ca3: x = 16'h1b2a; 14'h2ca4: x = 16'h1b29; 14'h2ca5: x = 16'h1b28; 14'h2ca6: x = 16'h1b27; 14'h2ca7: x = 16'h1b26; 14'h2ca8: x = 16'h1b26; 14'h2ca9: x = 16'h1b25; 14'h2caa: x = 16'h1b24; 14'h2cab: x = 16'h1b23; 14'h2cac: x = 16'h1b22; 14'h2cad: x = 16'h1b21; 14'h2cae: x = 16'h1b21; 14'h2caf: x = 16'h1b20; 14'h2cb0: x = 16'h1b1f; 14'h2cb1: x = 16'h1b1e; 14'h2cb2: x = 16'h1b1d; 14'h2cb3: x = 16'h1b1c; 14'h2cb4: x = 16'h1b1b; 14'h2cb5: x = 16'h1b1b; 14'h2cb6: x = 16'h1b1a; 14'h2cb7: x = 16'h1b19; 14'h2cb8: x = 16'h1b18; 14'h2cb9: x = 16'h1b17; 14'h2cba: x = 16'h1b16; 14'h2cbb: x = 16'h1b16; 14'h2cbc: x = 16'h1b15; 14'h2cbd: x = 16'h1b14; 14'h2cbe: x = 16'h1b13; 14'h2cbf: x = 16'h1b12; 14'h2cc0: x = 16'h1b11; 14'h2cc1: x = 16'h1b10; 14'h2cc2: x = 16'h1b10; 14'h2cc3: x = 16'h1b0f; 14'h2cc4: x = 16'h1b0e; 14'h2cc5: x = 16'h1b0d; 14'h2cc6: x = 16'h1b0c; 14'h2cc7: x = 16'h1b0b; 14'h2cc8: x = 16'h1b0b; 14'h2cc9: x = 16'h1b0a; 14'h2cca: x = 16'h1b09; 14'h2ccb: x = 16'h1b08; 14'h2ccc: x = 16'h1b07; 14'h2ccd: x = 16'h1b06; 14'h2cce: x = 16'h1b05; 14'h2ccf: x = 16'h1b05; 14'h2cd0: x = 16'h1b04; 14'h2cd1: x = 16'h1b03; 14'h2cd2: x = 16'h1b02; 14'h2cd3: x = 16'h1b01; 14'h2cd4: x = 16'h1b00; 14'h2cd5: x = 16'h1b00; 14'h2cd6: x = 16'h1aff; 14'h2cd7: x = 16'h1afe; 14'h2cd8: x = 16'h1afd; 14'h2cd9: x = 16'h1afc; 14'h2cda: x = 16'h1afb; 14'h2cdb: x = 16'h1afa; 14'h2cdc: x = 16'h1afa; 14'h2cdd: x = 16'h1af9; 14'h2cde: x = 16'h1af8; 14'h2cdf: x = 16'h1af7; 14'h2ce0: x = 16'h1af6; 14'h2ce1: x = 16'h1af5; 14'h2ce2: x = 16'h1af5; 14'h2ce3: x = 16'h1af4; 14'h2ce4: x = 16'h1af3; 14'h2ce5: x = 16'h1af2; 14'h2ce6: x = 16'h1af1; 14'h2ce7: x = 16'h1af0; 14'h2ce8: x = 16'h1aef; 14'h2ce9: x = 16'h1aef; 14'h2cea: x = 16'h1aee; 14'h2ceb: x = 16'h1aed; 14'h2cec: x = 16'h1aec; 14'h2ced: x = 16'h1aeb; 14'h2cee: x = 16'h1aea; 14'h2cef: x = 16'h1aea; 14'h2cf0: x = 16'h1ae9; 14'h2cf1: x = 16'h1ae8; 14'h2cf2: x = 16'h1ae7; 14'h2cf3: x = 16'h1ae6; 14'h2cf4: x = 16'h1ae5; 14'h2cf5: x = 16'h1ae4; 14'h2cf6: x = 16'h1ae4; 14'h2cf7: x = 16'h1ae3; 14'h2cf8: x = 16'h1ae2; 14'h2cf9: x = 16'h1ae1; 14'h2cfa: x = 16'h1ae0; 14'h2cfb: x = 16'h1adf; 14'h2cfc: x = 16'h1adf; 14'h2cfd: x = 16'h1ade; 14'h2cfe: x = 16'h1add; 14'h2cff: x = 16'h1adc; 14'h2d00: x = 16'h1adb; 14'h2d01: x = 16'h1ada; 14'h2d02: x = 16'h1ad9; 14'h2d03: x = 16'h1ad9; 14'h2d04: x = 16'h1ad8; 14'h2d05: x = 16'h1ad7; 14'h2d06: x = 16'h1ad6; 14'h2d07: x = 16'h1ad5; 14'h2d08: x = 16'h1ad4; 14'h2d09: x = 16'h1ad4; 14'h2d0a: x = 16'h1ad3; 14'h2d0b: x = 16'h1ad2; 14'h2d0c: x = 16'h1ad1; 14'h2d0d: x = 16'h1ad0; 14'h2d0e: x = 16'h1acf; 14'h2d0f: x = 16'h1ace; 14'h2d10: x = 16'h1ace; 14'h2d11: x = 16'h1acd; 14'h2d12: x = 16'h1acc; 14'h2d13: x = 16'h1acb; 14'h2d14: x = 16'h1aca; 14'h2d15: x = 16'h1ac9; 14'h2d16: x = 16'h1ac8; 14'h2d17: x = 16'h1ac8; 14'h2d18: x = 16'h1ac7; 14'h2d19: x = 16'h1ac6; 14'h2d1a: x = 16'h1ac5; 14'h2d1b: x = 16'h1ac4; 14'h2d1c: x = 16'h1ac3; 14'h2d1d: x = 16'h1ac3; 14'h2d1e: x = 16'h1ac2; 14'h2d1f: x = 16'h1ac1; 14'h2d20: x = 16'h1ac0; 14'h2d21: x = 16'h1abf; 14'h2d22: x = 16'h1abe; 14'h2d23: x = 16'h1abd; 14'h2d24: x = 16'h1abd; 14'h2d25: x = 16'h1abc; 14'h2d26: x = 16'h1abb; 14'h2d27: x = 16'h1aba; 14'h2d28: x = 16'h1ab9; 14'h2d29: x = 16'h1ab8; 14'h2d2a: x = 16'h1ab8; 14'h2d2b: x = 16'h1ab7; 14'h2d2c: x = 16'h1ab6; 14'h2d2d: x = 16'h1ab5; 14'h2d2e: x = 16'h1ab4; 14'h2d2f: x = 16'h1ab3; 14'h2d30: x = 16'h1ab2; 14'h2d31: x = 16'h1ab2; 14'h2d32: x = 16'h1ab1; 14'h2d33: x = 16'h1ab0; 14'h2d34: x = 16'h1aaf; 14'h2d35: x = 16'h1aae; 14'h2d36: x = 16'h1aad; 14'h2d37: x = 16'h1aac; 14'h2d38: x = 16'h1aac; 14'h2d39: x = 16'h1aab; 14'h2d3a: x = 16'h1aaa; 14'h2d3b: x = 16'h1aa9; 14'h2d3c: x = 16'h1aa8; 14'h2d3d: x = 16'h1aa7; 14'h2d3e: x = 16'h1aa7; 14'h2d3f: x = 16'h1aa6; 14'h2d40: x = 16'h1aa5; 14'h2d41: x = 16'h1aa4; 14'h2d42: x = 16'h1aa3; 14'h2d43: x = 16'h1aa2; 14'h2d44: x = 16'h1aa1; 14'h2d45: x = 16'h1aa1; 14'h2d46: x = 16'h1aa0; 14'h2d47: x = 16'h1a9f; 14'h2d48: x = 16'h1a9e; 14'h2d49: x = 16'h1a9d; 14'h2d4a: x = 16'h1a9c; 14'h2d4b: x = 16'h1a9b; 14'h2d4c: x = 16'h1a9b; 14'h2d4d: x = 16'h1a9a; 14'h2d4e: x = 16'h1a99; 14'h2d4f: x = 16'h1a98; 14'h2d50: x = 16'h1a97; 14'h2d51: x = 16'h1a96; 14'h2d52: x = 16'h1a96; 14'h2d53: x = 16'h1a95; 14'h2d54: x = 16'h1a94; 14'h2d55: x = 16'h1a93; 14'h2d56: x = 16'h1a92; 14'h2d57: x = 16'h1a91; 14'h2d58: x = 16'h1a90; 14'h2d59: x = 16'h1a90; 14'h2d5a: x = 16'h1a8f; 14'h2d5b: x = 16'h1a8e; 14'h2d5c: x = 16'h1a8d; 14'h2d5d: x = 16'h1a8c; 14'h2d5e: x = 16'h1a8b; 14'h2d5f: x = 16'h1a8a; 14'h2d60: x = 16'h1a8a; 14'h2d61: x = 16'h1a89; 14'h2d62: x = 16'h1a88; 14'h2d63: x = 16'h1a87; 14'h2d64: x = 16'h1a86; 14'h2d65: x = 16'h1a85; 14'h2d66: x = 16'h1a85; 14'h2d67: x = 16'h1a84; 14'h2d68: x = 16'h1a83; 14'h2d69: x = 16'h1a82; 14'h2d6a: x = 16'h1a81; 14'h2d6b: x = 16'h1a80; 14'h2d6c: x = 16'h1a7f; 14'h2d6d: x = 16'h1a7f; 14'h2d6e: x = 16'h1a7e; 14'h2d6f: x = 16'h1a7d; 14'h2d70: x = 16'h1a7c; 14'h2d71: x = 16'h1a7b; 14'h2d72: x = 16'h1a7a; 14'h2d73: x = 16'h1a79; 14'h2d74: x = 16'h1a79; 14'h2d75: x = 16'h1a78; 14'h2d76: x = 16'h1a77; 14'h2d77: x = 16'h1a76; 14'h2d78: x = 16'h1a75; 14'h2d79: x = 16'h1a74; 14'h2d7a: x = 16'h1a74; 14'h2d7b: x = 16'h1a73; 14'h2d7c: x = 16'h1a72; 14'h2d7d: x = 16'h1a71; 14'h2d7e: x = 16'h1a70; 14'h2d7f: x = 16'h1a6f; 14'h2d80: x = 16'h1a6e; 14'h2d81: x = 16'h1a6e; 14'h2d82: x = 16'h1a6d; 14'h2d83: x = 16'h1a6c; 14'h2d84: x = 16'h1a6b; 14'h2d85: x = 16'h1a6a; 14'h2d86: x = 16'h1a69; 14'h2d87: x = 16'h1a68; 14'h2d88: x = 16'h1a68; 14'h2d89: x = 16'h1a67; 14'h2d8a: x = 16'h1a66; 14'h2d8b: x = 16'h1a65; 14'h2d8c: x = 16'h1a64; 14'h2d8d: x = 16'h1a63; 14'h2d8e: x = 16'h1a62; 14'h2d8f: x = 16'h1a62; 14'h2d90: x = 16'h1a61; 14'h2d91: x = 16'h1a60; 14'h2d92: x = 16'h1a5f; 14'h2d93: x = 16'h1a5e; 14'h2d94: x = 16'h1a5d; 14'h2d95: x = 16'h1a5d; 14'h2d96: x = 16'h1a5c; 14'h2d97: x = 16'h1a5b; 14'h2d98: x = 16'h1a5a; 14'h2d99: x = 16'h1a59; 14'h2d9a: x = 16'h1a58; 14'h2d9b: x = 16'h1a57; 14'h2d9c: x = 16'h1a57; 14'h2d9d: x = 16'h1a56; 14'h2d9e: x = 16'h1a55; 14'h2d9f: x = 16'h1a54; 14'h2da0: x = 16'h1a53; 14'h2da1: x = 16'h1a52; 14'h2da2: x = 16'h1a51; 14'h2da3: x = 16'h1a51; 14'h2da4: x = 16'h1a50; 14'h2da5: x = 16'h1a4f; 14'h2da6: x = 16'h1a4e; 14'h2da7: x = 16'h1a4d; 14'h2da8: x = 16'h1a4c; 14'h2da9: x = 16'h1a4b; 14'h2daa: x = 16'h1a4b; 14'h2dab: x = 16'h1a4a; 14'h2dac: x = 16'h1a49; 14'h2dad: x = 16'h1a48; 14'h2dae: x = 16'h1a47; 14'h2daf: x = 16'h1a46; 14'h2db0: x = 16'h1a46; 14'h2db1: x = 16'h1a45; 14'h2db2: x = 16'h1a44; 14'h2db3: x = 16'h1a43; 14'h2db4: x = 16'h1a42; 14'h2db5: x = 16'h1a41; 14'h2db6: x = 16'h1a40; 14'h2db7: x = 16'h1a40; 14'h2db8: x = 16'h1a3f; 14'h2db9: x = 16'h1a3e; 14'h2dba: x = 16'h1a3d; 14'h2dbb: x = 16'h1a3c; 14'h2dbc: x = 16'h1a3b; 14'h2dbd: x = 16'h1a3a; 14'h2dbe: x = 16'h1a3a; 14'h2dbf: x = 16'h1a39; 14'h2dc0: x = 16'h1a38; 14'h2dc1: x = 16'h1a37; 14'h2dc2: x = 16'h1a36; 14'h2dc3: x = 16'h1a35; 14'h2dc4: x = 16'h1a34; 14'h2dc5: x = 16'h1a34; 14'h2dc6: x = 16'h1a33; 14'h2dc7: x = 16'h1a32; 14'h2dc8: x = 16'h1a31; 14'h2dc9: x = 16'h1a30; 14'h2dca: x = 16'h1a2f; 14'h2dcb: x = 16'h1a2e; 14'h2dcc: x = 16'h1a2e; 14'h2dcd: x = 16'h1a2d; 14'h2dce: x = 16'h1a2c; 14'h2dcf: x = 16'h1a2b; 14'h2dd0: x = 16'h1a2a; 14'h2dd1: x = 16'h1a29; 14'h2dd2: x = 16'h1a28; 14'h2dd3: x = 16'h1a28; 14'h2dd4: x = 16'h1a27; 14'h2dd5: x = 16'h1a26; 14'h2dd6: x = 16'h1a25; 14'h2dd7: x = 16'h1a24; 14'h2dd8: x = 16'h1a23; 14'h2dd9: x = 16'h1a23; 14'h2dda: x = 16'h1a22; 14'h2ddb: x = 16'h1a21; 14'h2ddc: x = 16'h1a20; 14'h2ddd: x = 16'h1a1f; 14'h2dde: x = 16'h1a1e; 14'h2ddf: x = 16'h1a1d; 14'h2de0: x = 16'h1a1d; 14'h2de1: x = 16'h1a1c; 14'h2de2: x = 16'h1a1b; 14'h2de3: x = 16'h1a1a; 14'h2de4: x = 16'h1a19; 14'h2de5: x = 16'h1a18; 14'h2de6: x = 16'h1a17; 14'h2de7: x = 16'h1a17; 14'h2de8: x = 16'h1a16; 14'h2de9: x = 16'h1a15; 14'h2dea: x = 16'h1a14; 14'h2deb: x = 16'h1a13; 14'h2dec: x = 16'h1a12; 14'h2ded: x = 16'h1a11; 14'h2dee: x = 16'h1a11; 14'h2def: x = 16'h1a10; 14'h2df0: x = 16'h1a0f; 14'h2df1: x = 16'h1a0e; 14'h2df2: x = 16'h1a0d; 14'h2df3: x = 16'h1a0c; 14'h2df4: x = 16'h1a0b; 14'h2df5: x = 16'h1a0b; 14'h2df6: x = 16'h1a0a; 14'h2df7: x = 16'h1a09; 14'h2df8: x = 16'h1a08; 14'h2df9: x = 16'h1a07; 14'h2dfa: x = 16'h1a06; 14'h2dfb: x = 16'h1a05; 14'h2dfc: x = 16'h1a05; 14'h2dfd: x = 16'h1a04; 14'h2dfe: x = 16'h1a03; 14'h2dff: x = 16'h1a02; 14'h2e00: x = 16'h1a01; 14'h2e01: x = 16'h1a00; 14'h2e02: x = 16'h19ff; 14'h2e03: x = 16'h19ff; 14'h2e04: x = 16'h19fe; 14'h2e05: x = 16'h19fd; 14'h2e06: x = 16'h19fc; 14'h2e07: x = 16'h19fb; 14'h2e08: x = 16'h19fa; 14'h2e09: x = 16'h19f9; 14'h2e0a: x = 16'h19f9; 14'h2e0b: x = 16'h19f8; 14'h2e0c: x = 16'h19f7; 14'h2e0d: x = 16'h19f6; 14'h2e0e: x = 16'h19f5; 14'h2e0f: x = 16'h19f4; 14'h2e10: x = 16'h19f3; 14'h2e11: x = 16'h19f3; 14'h2e12: x = 16'h19f2; 14'h2e13: x = 16'h19f1; 14'h2e14: x = 16'h19f0; 14'h2e15: x = 16'h19ef; 14'h2e16: x = 16'h19ee; 14'h2e17: x = 16'h19ed; 14'h2e18: x = 16'h19ed; 14'h2e19: x = 16'h19ec; 14'h2e1a: x = 16'h19eb; 14'h2e1b: x = 16'h19ea; 14'h2e1c: x = 16'h19e9; 14'h2e1d: x = 16'h19e8; 14'h2e1e: x = 16'h19e7; 14'h2e1f: x = 16'h19e7; 14'h2e20: x = 16'h19e6; 14'h2e21: x = 16'h19e5; 14'h2e22: x = 16'h19e4; 14'h2e23: x = 16'h19e3; 14'h2e24: x = 16'h19e2; 14'h2e25: x = 16'h19e1; 14'h2e26: x = 16'h19e1; 14'h2e27: x = 16'h19e0; 14'h2e28: x = 16'h19df; 14'h2e29: x = 16'h19de; 14'h2e2a: x = 16'h19dd; 14'h2e2b: x = 16'h19dc; 14'h2e2c: x = 16'h19db; 14'h2e2d: x = 16'h19db; 14'h2e2e: x = 16'h19da; 14'h2e2f: x = 16'h19d9; 14'h2e30: x = 16'h19d8; 14'h2e31: x = 16'h19d7; 14'h2e32: x = 16'h19d6; 14'h2e33: x = 16'h19d5; 14'h2e34: x = 16'h19d5; 14'h2e35: x = 16'h19d4; 14'h2e36: x = 16'h19d3; 14'h2e37: x = 16'h19d2; 14'h2e38: x = 16'h19d1; 14'h2e39: x = 16'h19d0; 14'h2e3a: x = 16'h19cf; 14'h2e3b: x = 16'h19cf; 14'h2e3c: x = 16'h19ce; 14'h2e3d: x = 16'h19cd; 14'h2e3e: x = 16'h19cc; 14'h2e3f: x = 16'h19cb; 14'h2e40: x = 16'h19ca; 14'h2e41: x = 16'h19c9; 14'h2e42: x = 16'h19c9; 14'h2e43: x = 16'h19c8; 14'h2e44: x = 16'h19c7; 14'h2e45: x = 16'h19c6; 14'h2e46: x = 16'h19c5; 14'h2e47: x = 16'h19c4; 14'h2e48: x = 16'h19c3; 14'h2e49: x = 16'h19c3; 14'h2e4a: x = 16'h19c2; 14'h2e4b: x = 16'h19c1; 14'h2e4c: x = 16'h19c0; 14'h2e4d: x = 16'h19bf; 14'h2e4e: x = 16'h19be; 14'h2e4f: x = 16'h19bd; 14'h2e50: x = 16'h19bd; 14'h2e51: x = 16'h19bc; 14'h2e52: x = 16'h19bb; 14'h2e53: x = 16'h19ba; 14'h2e54: x = 16'h19b9; 14'h2e55: x = 16'h19b8; 14'h2e56: x = 16'h19b7; 14'h2e57: x = 16'h19b7; 14'h2e58: x = 16'h19b6; 14'h2e59: x = 16'h19b5; 14'h2e5a: x = 16'h19b4; 14'h2e5b: x = 16'h19b3; 14'h2e5c: x = 16'h19b2; 14'h2e5d: x = 16'h19b1; 14'h2e5e: x = 16'h19b1; 14'h2e5f: x = 16'h19b0; 14'h2e60: x = 16'h19af; 14'h2e61: x = 16'h19ae; 14'h2e62: x = 16'h19ad; 14'h2e63: x = 16'h19ac; 14'h2e64: x = 16'h19ab; 14'h2e65: x = 16'h19ab; 14'h2e66: x = 16'h19aa; 14'h2e67: x = 16'h19a9; 14'h2e68: x = 16'h19a8; 14'h2e69: x = 16'h19a7; 14'h2e6a: x = 16'h19a6; 14'h2e6b: x = 16'h19a5; 14'h2e6c: x = 16'h19a4; 14'h2e6d: x = 16'h19a4; 14'h2e6e: x = 16'h19a3; 14'h2e6f: x = 16'h19a2; 14'h2e70: x = 16'h19a1; 14'h2e71: x = 16'h19a0; 14'h2e72: x = 16'h199f; 14'h2e73: x = 16'h199e; 14'h2e74: x = 16'h199e; 14'h2e75: x = 16'h199d; 14'h2e76: x = 16'h199c; 14'h2e77: x = 16'h199b; 14'h2e78: x = 16'h199a; 14'h2e79: x = 16'h1999; 14'h2e7a: x = 16'h1998; 14'h2e7b: x = 16'h1998; 14'h2e7c: x = 16'h1997; 14'h2e7d: x = 16'h1996; 14'h2e7e: x = 16'h1995; 14'h2e7f: x = 16'h1994; 14'h2e80: x = 16'h1993; 14'h2e81: x = 16'h1992; 14'h2e82: x = 16'h1992; 14'h2e83: x = 16'h1991; 14'h2e84: x = 16'h1990; 14'h2e85: x = 16'h198f; 14'h2e86: x = 16'h198e; 14'h2e87: x = 16'h198d; 14'h2e88: x = 16'h198c; 14'h2e89: x = 16'h198c; 14'h2e8a: x = 16'h198b; 14'h2e8b: x = 16'h198a; 14'h2e8c: x = 16'h1989; 14'h2e8d: x = 16'h1988; 14'h2e8e: x = 16'h1987; 14'h2e8f: x = 16'h1986; 14'h2e90: x = 16'h1985; 14'h2e91: x = 16'h1985; 14'h2e92: x = 16'h1984; 14'h2e93: x = 16'h1983; 14'h2e94: x = 16'h1982; 14'h2e95: x = 16'h1981; 14'h2e96: x = 16'h1980; 14'h2e97: x = 16'h197f; 14'h2e98: x = 16'h197f; 14'h2e99: x = 16'h197e; 14'h2e9a: x = 16'h197d; 14'h2e9b: x = 16'h197c; 14'h2e9c: x = 16'h197b; 14'h2e9d: x = 16'h197a; 14'h2e9e: x = 16'h1979; 14'h2e9f: x = 16'h1979; 14'h2ea0: x = 16'h1978; 14'h2ea1: x = 16'h1977; 14'h2ea2: x = 16'h1976; 14'h2ea3: x = 16'h1975; 14'h2ea4: x = 16'h1974; 14'h2ea5: x = 16'h1973; 14'h2ea6: x = 16'h1973; 14'h2ea7: x = 16'h1972; 14'h2ea8: x = 16'h1971; 14'h2ea9: x = 16'h1970; 14'h2eaa: x = 16'h196f; 14'h2eab: x = 16'h196e; 14'h2eac: x = 16'h196d; 14'h2ead: x = 16'h196c; 14'h2eae: x = 16'h196c; 14'h2eaf: x = 16'h196b; 14'h2eb0: x = 16'h196a; 14'h2eb1: x = 16'h1969; 14'h2eb2: x = 16'h1968; 14'h2eb3: x = 16'h1967; 14'h2eb4: x = 16'h1966; 14'h2eb5: x = 16'h1966; 14'h2eb6: x = 16'h1965; 14'h2eb7: x = 16'h1964; 14'h2eb8: x = 16'h1963; 14'h2eb9: x = 16'h1962; 14'h2eba: x = 16'h1961; 14'h2ebb: x = 16'h1960; 14'h2ebc: x = 16'h1960; 14'h2ebd: x = 16'h195f; 14'h2ebe: x = 16'h195e; 14'h2ebf: x = 16'h195d; 14'h2ec0: x = 16'h195c; 14'h2ec1: x = 16'h195b; 14'h2ec2: x = 16'h195a; 14'h2ec3: x = 16'h1959; 14'h2ec4: x = 16'h1959; 14'h2ec5: x = 16'h1958; 14'h2ec6: x = 16'h1957; 14'h2ec7: x = 16'h1956; 14'h2ec8: x = 16'h1955; 14'h2ec9: x = 16'h1954; 14'h2eca: x = 16'h1953; 14'h2ecb: x = 16'h1953; 14'h2ecc: x = 16'h1952; 14'h2ecd: x = 16'h1951; 14'h2ece: x = 16'h1950; 14'h2ecf: x = 16'h194f; 14'h2ed0: x = 16'h194e; 14'h2ed1: x = 16'h194d; 14'h2ed2: x = 16'h194d; 14'h2ed3: x = 16'h194c; 14'h2ed4: x = 16'h194b; 14'h2ed5: x = 16'h194a; 14'h2ed6: x = 16'h1949; 14'h2ed7: x = 16'h1948; 14'h2ed8: x = 16'h1947; 14'h2ed9: x = 16'h1946; 14'h2eda: x = 16'h1946; 14'h2edb: x = 16'h1945; 14'h2edc: x = 16'h1944; 14'h2edd: x = 16'h1943; 14'h2ede: x = 16'h1942; 14'h2edf: x = 16'h1941; 14'h2ee0: x = 16'h1940; 14'h2ee1: x = 16'h1940; 14'h2ee2: x = 16'h193f; 14'h2ee3: x = 16'h193e; 14'h2ee4: x = 16'h193d; 14'h2ee5: x = 16'h193c; 14'h2ee6: x = 16'h193b; 14'h2ee7: x = 16'h193a; 14'h2ee8: x = 16'h1939; 14'h2ee9: x = 16'h1939; 14'h2eea: x = 16'h1938; 14'h2eeb: x = 16'h1937; 14'h2eec: x = 16'h1936; 14'h2eed: x = 16'h1935; 14'h2eee: x = 16'h1934; 14'h2eef: x = 16'h1933; 14'h2ef0: x = 16'h1933; 14'h2ef1: x = 16'h1932; 14'h2ef2: x = 16'h1931; 14'h2ef3: x = 16'h1930; 14'h2ef4: x = 16'h192f; 14'h2ef5: x = 16'h192e; 14'h2ef6: x = 16'h192d; 14'h2ef7: x = 16'h192d; 14'h2ef8: x = 16'h192c; 14'h2ef9: x = 16'h192b; 14'h2efa: x = 16'h192a; 14'h2efb: x = 16'h1929; 14'h2efc: x = 16'h1928; 14'h2efd: x = 16'h1927; 14'h2efe: x = 16'h1926; 14'h2eff: x = 16'h1926; 14'h2f00: x = 16'h1925; 14'h2f01: x = 16'h1924; 14'h2f02: x = 16'h1923; 14'h2f03: x = 16'h1922; 14'h2f04: x = 16'h1921; 14'h2f05: x = 16'h1920; 14'h2f06: x = 16'h1920; 14'h2f07: x = 16'h191f; 14'h2f08: x = 16'h191e; 14'h2f09: x = 16'h191d; 14'h2f0a: x = 16'h191c; 14'h2f0b: x = 16'h191b; 14'h2f0c: x = 16'h191a; 14'h2f0d: x = 16'h1919; 14'h2f0e: x = 16'h1919; 14'h2f0f: x = 16'h1918; 14'h2f10: x = 16'h1917; 14'h2f11: x = 16'h1916; 14'h2f12: x = 16'h1915; 14'h2f13: x = 16'h1914; 14'h2f14: x = 16'h1913; 14'h2f15: x = 16'h1913; 14'h2f16: x = 16'h1912; 14'h2f17: x = 16'h1911; 14'h2f18: x = 16'h1910; 14'h2f19: x = 16'h190f; 14'h2f1a: x = 16'h190e; 14'h2f1b: x = 16'h190d; 14'h2f1c: x = 16'h190c; 14'h2f1d: x = 16'h190c; 14'h2f1e: x = 16'h190b; 14'h2f1f: x = 16'h190a; 14'h2f20: x = 16'h1909; 14'h2f21: x = 16'h1908; 14'h2f22: x = 16'h1907; 14'h2f23: x = 16'h1906; 14'h2f24: x = 16'h1905; 14'h2f25: x = 16'h1905; 14'h2f26: x = 16'h1904; 14'h2f27: x = 16'h1903; 14'h2f28: x = 16'h1902; 14'h2f29: x = 16'h1901; 14'h2f2a: x = 16'h1900; 14'h2f2b: x = 16'h18ff; 14'h2f2c: x = 16'h18ff; 14'h2f2d: x = 16'h18fe; 14'h2f2e: x = 16'h18fd; 14'h2f2f: x = 16'h18fc; 14'h2f30: x = 16'h18fb; 14'h2f31: x = 16'h18fa; 14'h2f32: x = 16'h18f9; 14'h2f33: x = 16'h18f8; 14'h2f34: x = 16'h18f8; 14'h2f35: x = 16'h18f7; 14'h2f36: x = 16'h18f6; 14'h2f37: x = 16'h18f5; 14'h2f38: x = 16'h18f4; 14'h2f39: x = 16'h18f3; 14'h2f3a: x = 16'h18f2; 14'h2f3b: x = 16'h18f2; 14'h2f3c: x = 16'h18f1; 14'h2f3d: x = 16'h18f0; 14'h2f3e: x = 16'h18ef; 14'h2f3f: x = 16'h18ee; 14'h2f40: x = 16'h18ed; 14'h2f41: x = 16'h18ec; 14'h2f42: x = 16'h18eb; 14'h2f43: x = 16'h18eb; 14'h2f44: x = 16'h18ea; 14'h2f45: x = 16'h18e9; 14'h2f46: x = 16'h18e8; 14'h2f47: x = 16'h18e7; 14'h2f48: x = 16'h18e6; 14'h2f49: x = 16'h18e5; 14'h2f4a: x = 16'h18e4; 14'h2f4b: x = 16'h18e4; 14'h2f4c: x = 16'h18e3; 14'h2f4d: x = 16'h18e2; 14'h2f4e: x = 16'h18e1; 14'h2f4f: x = 16'h18e0; 14'h2f50: x = 16'h18df; 14'h2f51: x = 16'h18de; 14'h2f52: x = 16'h18de; 14'h2f53: x = 16'h18dd; 14'h2f54: x = 16'h18dc; 14'h2f55: x = 16'h18db; 14'h2f56: x = 16'h18da; 14'h2f57: x = 16'h18d9; 14'h2f58: x = 16'h18d8; 14'h2f59: x = 16'h18d7; 14'h2f5a: x = 16'h18d7; 14'h2f5b: x = 16'h18d6; 14'h2f5c: x = 16'h18d5; 14'h2f5d: x = 16'h18d4; 14'h2f5e: x = 16'h18d3; 14'h2f5f: x = 16'h18d2; 14'h2f60: x = 16'h18d1; 14'h2f61: x = 16'h18d0; 14'h2f62: x = 16'h18d0; 14'h2f63: x = 16'h18cf; 14'h2f64: x = 16'h18ce; 14'h2f65: x = 16'h18cd; 14'h2f66: x = 16'h18cc; 14'h2f67: x = 16'h18cb; 14'h2f68: x = 16'h18ca; 14'h2f69: x = 16'h18c9; 14'h2f6a: x = 16'h18c9; 14'h2f6b: x = 16'h18c8; 14'h2f6c: x = 16'h18c7; 14'h2f6d: x = 16'h18c6; 14'h2f6e: x = 16'h18c5; 14'h2f6f: x = 16'h18c4; 14'h2f70: x = 16'h18c3; 14'h2f71: x = 16'h18c3; 14'h2f72: x = 16'h18c2; 14'h2f73: x = 16'h18c1; 14'h2f74: x = 16'h18c0; 14'h2f75: x = 16'h18bf; 14'h2f76: x = 16'h18be; 14'h2f77: x = 16'h18bd; 14'h2f78: x = 16'h18bc; 14'h2f79: x = 16'h18bc; 14'h2f7a: x = 16'h18bb; 14'h2f7b: x = 16'h18ba; 14'h2f7c: x = 16'h18b9; 14'h2f7d: x = 16'h18b8; 14'h2f7e: x = 16'h18b7; 14'h2f7f: x = 16'h18b6; 14'h2f80: x = 16'h18b5; 14'h2f81: x = 16'h18b5; 14'h2f82: x = 16'h18b4; 14'h2f83: x = 16'h18b3; 14'h2f84: x = 16'h18b2; 14'h2f85: x = 16'h18b1; 14'h2f86: x = 16'h18b0; 14'h2f87: x = 16'h18af; 14'h2f88: x = 16'h18ae; 14'h2f89: x = 16'h18ae; 14'h2f8a: x = 16'h18ad; 14'h2f8b: x = 16'h18ac; 14'h2f8c: x = 16'h18ab; 14'h2f8d: x = 16'h18aa; 14'h2f8e: x = 16'h18a9; 14'h2f8f: x = 16'h18a8; 14'h2f90: x = 16'h18a7; 14'h2f91: x = 16'h18a7; 14'h2f92: x = 16'h18a6; 14'h2f93: x = 16'h18a5; 14'h2f94: x = 16'h18a4; 14'h2f95: x = 16'h18a3; 14'h2f96: x = 16'h18a2; 14'h2f97: x = 16'h18a1; 14'h2f98: x = 16'h18a0; 14'h2f99: x = 16'h18a0; 14'h2f9a: x = 16'h189f; 14'h2f9b: x = 16'h189e; 14'h2f9c: x = 16'h189d; 14'h2f9d: x = 16'h189c; 14'h2f9e: x = 16'h189b; 14'h2f9f: x = 16'h189a; 14'h2fa0: x = 16'h1899; 14'h2fa1: x = 16'h1899; 14'h2fa2: x = 16'h1898; 14'h2fa3: x = 16'h1897; 14'h2fa4: x = 16'h1896; 14'h2fa5: x = 16'h1895; 14'h2fa6: x = 16'h1894; 14'h2fa7: x = 16'h1893; 14'h2fa8: x = 16'h1893; 14'h2fa9: x = 16'h1892; 14'h2faa: x = 16'h1891; 14'h2fab: x = 16'h1890; 14'h2fac: x = 16'h188f; 14'h2fad: x = 16'h188e; 14'h2fae: x = 16'h188d; 14'h2faf: x = 16'h188c; 14'h2fb0: x = 16'h188c; 14'h2fb1: x = 16'h188b; 14'h2fb2: x = 16'h188a; 14'h2fb3: x = 16'h1889; 14'h2fb4: x = 16'h1888; 14'h2fb5: x = 16'h1887; 14'h2fb6: x = 16'h1886; 14'h2fb7: x = 16'h1885; 14'h2fb8: x = 16'h1885; 14'h2fb9: x = 16'h1884; 14'h2fba: x = 16'h1883; 14'h2fbb: x = 16'h1882; 14'h2fbc: x = 16'h1881; 14'h2fbd: x = 16'h1880; 14'h2fbe: x = 16'h187f; 14'h2fbf: x = 16'h187e; 14'h2fc0: x = 16'h187e; 14'h2fc1: x = 16'h187d; 14'h2fc2: x = 16'h187c; 14'h2fc3: x = 16'h187b; 14'h2fc4: x = 16'h187a; 14'h2fc5: x = 16'h1879; 14'h2fc6: x = 16'h1878; 14'h2fc7: x = 16'h1877; 14'h2fc8: x = 16'h1876; 14'h2fc9: x = 16'h1876; 14'h2fca: x = 16'h1875; 14'h2fcb: x = 16'h1874; 14'h2fcc: x = 16'h1873; 14'h2fcd: x = 16'h1872; 14'h2fce: x = 16'h1871; 14'h2fcf: x = 16'h1870; 14'h2fd0: x = 16'h186f; 14'h2fd1: x = 16'h186f; 14'h2fd2: x = 16'h186e; 14'h2fd3: x = 16'h186d; 14'h2fd4: x = 16'h186c; 14'h2fd5: x = 16'h186b; 14'h2fd6: x = 16'h186a; 14'h2fd7: x = 16'h1869; 14'h2fd8: x = 16'h1868; 14'h2fd9: x = 16'h1868; 14'h2fda: x = 16'h1867; 14'h2fdb: x = 16'h1866; 14'h2fdc: x = 16'h1865; 14'h2fdd: x = 16'h1864; 14'h2fde: x = 16'h1863; 14'h2fdf: x = 16'h1862; 14'h2fe0: x = 16'h1861; 14'h2fe1: x = 16'h1861; 14'h2fe2: x = 16'h1860; 14'h2fe3: x = 16'h185f; 14'h2fe4: x = 16'h185e; 14'h2fe5: x = 16'h185d; 14'h2fe6: x = 16'h185c; 14'h2fe7: x = 16'h185b; 14'h2fe8: x = 16'h185a; 14'h2fe9: x = 16'h185a; 14'h2fea: x = 16'h1859; 14'h2feb: x = 16'h1858; 14'h2fec: x = 16'h1857; 14'h2fed: x = 16'h1856; 14'h2fee: x = 16'h1855; 14'h2fef: x = 16'h1854; 14'h2ff0: x = 16'h1853; 14'h2ff1: x = 16'h1853; 14'h2ff2: x = 16'h1852; 14'h2ff3: x = 16'h1851; 14'h2ff4: x = 16'h1850; 14'h2ff5: x = 16'h184f; 14'h2ff6: x = 16'h184e; 14'h2ff7: x = 16'h184d; 14'h2ff8: x = 16'h184c; 14'h2ff9: x = 16'h184c; 14'h2ffa: x = 16'h184b; 14'h2ffb: x = 16'h184a; 14'h2ffc: x = 16'h1849; 14'h2ffd: x = 16'h1848; 14'h2ffe: x = 16'h1847; 14'h2fff: x = 16'h1846; 14'h3000: x = 16'h1845; 14'h3001: x = 16'h1844; 14'h3002: x = 16'h1844; 14'h3003: x = 16'h1843; 14'h3004: x = 16'h1842; 14'h3005: x = 16'h1841; 14'h3006: x = 16'h1840; 14'h3007: x = 16'h183f; 14'h3008: x = 16'h183e; 14'h3009: x = 16'h183d; 14'h300a: x = 16'h183d; 14'h300b: x = 16'h183c; 14'h300c: x = 16'h183b; 14'h300d: x = 16'h183a; 14'h300e: x = 16'h1839; 14'h300f: x = 16'h1838; 14'h3010: x = 16'h1837; 14'h3011: x = 16'h1836; 14'h3012: x = 16'h1836; 14'h3013: x = 16'h1835; 14'h3014: x = 16'h1834; 14'h3015: x = 16'h1833; 14'h3016: x = 16'h1832; 14'h3017: x = 16'h1831; 14'h3018: x = 16'h1830; 14'h3019: x = 16'h182f; 14'h301a: x = 16'h182e; 14'h301b: x = 16'h182e; 14'h301c: x = 16'h182d; 14'h301d: x = 16'h182c; 14'h301e: x = 16'h182b; 14'h301f: x = 16'h182a; 14'h3020: x = 16'h1829; 14'h3021: x = 16'h1828; 14'h3022: x = 16'h1827; 14'h3023: x = 16'h1827; 14'h3024: x = 16'h1826; 14'h3025: x = 16'h1825; 14'h3026: x = 16'h1824; 14'h3027: x = 16'h1823; 14'h3028: x = 16'h1822; 14'h3029: x = 16'h1821; 14'h302a: x = 16'h1820; 14'h302b: x = 16'h1820; 14'h302c: x = 16'h181f; 14'h302d: x = 16'h181e; 14'h302e: x = 16'h181d; 14'h302f: x = 16'h181c; 14'h3030: x = 16'h181b; 14'h3031: x = 16'h181a; 14'h3032: x = 16'h1819; 14'h3033: x = 16'h1818; 14'h3034: x = 16'h1818; 14'h3035: x = 16'h1817; 14'h3036: x = 16'h1816; 14'h3037: x = 16'h1815; 14'h3038: x = 16'h1814; 14'h3039: x = 16'h1813; 14'h303a: x = 16'h1812; 14'h303b: x = 16'h1811; 14'h303c: x = 16'h1811; 14'h303d: x = 16'h1810; 14'h303e: x = 16'h180f; 14'h303f: x = 16'h180e; 14'h3040: x = 16'h180d; 14'h3041: x = 16'h180c; 14'h3042: x = 16'h180b; 14'h3043: x = 16'h180a; 14'h3044: x = 16'h1809; 14'h3045: x = 16'h1809; 14'h3046: x = 16'h1808; 14'h3047: x = 16'h1807; 14'h3048: x = 16'h1806; 14'h3049: x = 16'h1805; 14'h304a: x = 16'h1804; 14'h304b: x = 16'h1803; 14'h304c: x = 16'h1802; 14'h304d: x = 16'h1802; 14'h304e: x = 16'h1801; 14'h304f: x = 16'h1800; 14'h3050: x = 16'h17ff; 14'h3051: x = 16'h17fe; 14'h3052: x = 16'h17fd; 14'h3053: x = 16'h17fc; 14'h3054: x = 16'h17fb; 14'h3055: x = 16'h17fa; 14'h3056: x = 16'h17fa; 14'h3057: x = 16'h17f9; 14'h3058: x = 16'h17f8; 14'h3059: x = 16'h17f7; 14'h305a: x = 16'h17f6; 14'h305b: x = 16'h17f5; 14'h305c: x = 16'h17f4; 14'h305d: x = 16'h17f3; 14'h305e: x = 16'h17f3; 14'h305f: x = 16'h17f2; 14'h3060: x = 16'h17f1; 14'h3061: x = 16'h17f0; 14'h3062: x = 16'h17ef; 14'h3063: x = 16'h17ee; 14'h3064: x = 16'h17ed; 14'h3065: x = 16'h17ec; 14'h3066: x = 16'h17eb; 14'h3067: x = 16'h17eb; 14'h3068: x = 16'h17ea; 14'h3069: x = 16'h17e9; 14'h306a: x = 16'h17e8; 14'h306b: x = 16'h17e7; 14'h306c: x = 16'h17e6; 14'h306d: x = 16'h17e5; 14'h306e: x = 16'h17e4; 14'h306f: x = 16'h17e3; 14'h3070: x = 16'h17e3; 14'h3071: x = 16'h17e2; 14'h3072: x = 16'h17e1; 14'h3073: x = 16'h17e0; 14'h3074: x = 16'h17df; 14'h3075: x = 16'h17de; 14'h3076: x = 16'h17dd; 14'h3077: x = 16'h17dc; 14'h3078: x = 16'h17dc; 14'h3079: x = 16'h17db; 14'h307a: x = 16'h17da; 14'h307b: x = 16'h17d9; 14'h307c: x = 16'h17d8; 14'h307d: x = 16'h17d7; 14'h307e: x = 16'h17d6; 14'h307f: x = 16'h17d5; 14'h3080: x = 16'h17d4; 14'h3081: x = 16'h17d4; 14'h3082: x = 16'h17d3; 14'h3083: x = 16'h17d2; 14'h3084: x = 16'h17d1; 14'h3085: x = 16'h17d0; 14'h3086: x = 16'h17cf; 14'h3087: x = 16'h17ce; 14'h3088: x = 16'h17cd; 14'h3089: x = 16'h17cc; 14'h308a: x = 16'h17cc; 14'h308b: x = 16'h17cb; 14'h308c: x = 16'h17ca; 14'h308d: x = 16'h17c9; 14'h308e: x = 16'h17c8; 14'h308f: x = 16'h17c7; 14'h3090: x = 16'h17c6; 14'h3091: x = 16'h17c5; 14'h3092: x = 16'h17c4; 14'h3093: x = 16'h17c4; 14'h3094: x = 16'h17c3; 14'h3095: x = 16'h17c2; 14'h3096: x = 16'h17c1; 14'h3097: x = 16'h17c0; 14'h3098: x = 16'h17bf; 14'h3099: x = 16'h17be; 14'h309a: x = 16'h17bd; 14'h309b: x = 16'h17bc; 14'h309c: x = 16'h17bc; 14'h309d: x = 16'h17bb; 14'h309e: x = 16'h17ba; 14'h309f: x = 16'h17b9; 14'h30a0: x = 16'h17b8; 14'h30a1: x = 16'h17b7; 14'h30a2: x = 16'h17b6; 14'h30a3: x = 16'h17b5; 14'h30a4: x = 16'h17b4; 14'h30a5: x = 16'h17b4; 14'h30a6: x = 16'h17b3; 14'h30a7: x = 16'h17b2; 14'h30a8: x = 16'h17b1; 14'h30a9: x = 16'h17b0; 14'h30aa: x = 16'h17af; 14'h30ab: x = 16'h17ae; 14'h30ac: x = 16'h17ad; 14'h30ad: x = 16'h17ac; 14'h30ae: x = 16'h17ac; 14'h30af: x = 16'h17ab; 14'h30b0: x = 16'h17aa; 14'h30b1: x = 16'h17a9; 14'h30b2: x = 16'h17a8; 14'h30b3: x = 16'h17a7; 14'h30b4: x = 16'h17a6; 14'h30b5: x = 16'h17a5; 14'h30b6: x = 16'h17a4; 14'h30b7: x = 16'h17a4; 14'h30b8: x = 16'h17a3; 14'h30b9: x = 16'h17a2; 14'h30ba: x = 16'h17a1; 14'h30bb: x = 16'h17a0; 14'h30bc: x = 16'h179f; 14'h30bd: x = 16'h179e; 14'h30be: x = 16'h179d; 14'h30bf: x = 16'h179c; 14'h30c0: x = 16'h179c; 14'h30c1: x = 16'h179b; 14'h30c2: x = 16'h179a; 14'h30c3: x = 16'h1799; 14'h30c4: x = 16'h1798; 14'h30c5: x = 16'h1797; 14'h30c6: x = 16'h1796; 14'h30c7: x = 16'h1795; 14'h30c8: x = 16'h1794; 14'h30c9: x = 16'h1794; 14'h30ca: x = 16'h1793; 14'h30cb: x = 16'h1792; 14'h30cc: x = 16'h1791; 14'h30cd: x = 16'h1790; 14'h30ce: x = 16'h178f; 14'h30cf: x = 16'h178e; 14'h30d0: x = 16'h178d; 14'h30d1: x = 16'h178c; 14'h30d2: x = 16'h178c; 14'h30d3: x = 16'h178b; 14'h30d4: x = 16'h178a; 14'h30d5: x = 16'h1789; 14'h30d6: x = 16'h1788; 14'h30d7: x = 16'h1787; 14'h30d8: x = 16'h1786; 14'h30d9: x = 16'h1785; 14'h30da: x = 16'h1784; 14'h30db: x = 16'h1784; 14'h30dc: x = 16'h1783; 14'h30dd: x = 16'h1782; 14'h30de: x = 16'h1781; 14'h30df: x = 16'h1780; 14'h30e0: x = 16'h177f; 14'h30e1: x = 16'h177e; 14'h30e2: x = 16'h177d; 14'h30e3: x = 16'h177c; 14'h30e4: x = 16'h177c; 14'h30e5: x = 16'h177b; 14'h30e6: x = 16'h177a; 14'h30e7: x = 16'h1779; 14'h30e8: x = 16'h1778; 14'h30e9: x = 16'h1777; 14'h30ea: x = 16'h1776; 14'h30eb: x = 16'h1775; 14'h30ec: x = 16'h1774; 14'h30ed: x = 16'h1773; 14'h30ee: x = 16'h1773; 14'h30ef: x = 16'h1772; 14'h30f0: x = 16'h1771; 14'h30f1: x = 16'h1770; 14'h30f2: x = 16'h176f; 14'h30f3: x = 16'h176e; 14'h30f4: x = 16'h176d; 14'h30f5: x = 16'h176c; 14'h30f6: x = 16'h176b; 14'h30f7: x = 16'h176b; 14'h30f8: x = 16'h176a; 14'h30f9: x = 16'h1769; 14'h30fa: x = 16'h1768; 14'h30fb: x = 16'h1767; 14'h30fc: x = 16'h1766; 14'h30fd: x = 16'h1765; 14'h30fe: x = 16'h1764; 14'h30ff: x = 16'h1763; 14'h3100: x = 16'h1763; 14'h3101: x = 16'h1762; 14'h3102: x = 16'h1761; 14'h3103: x = 16'h1760; 14'h3104: x = 16'h175f; 14'h3105: x = 16'h175e; 14'h3106: x = 16'h175d; 14'h3107: x = 16'h175c; 14'h3108: x = 16'h175b; 14'h3109: x = 16'h175a; 14'h310a: x = 16'h175a; 14'h310b: x = 16'h1759; 14'h310c: x = 16'h1758; 14'h310d: x = 16'h1757; 14'h310e: x = 16'h1756; 14'h310f: x = 16'h1755; 14'h3110: x = 16'h1754; 14'h3111: x = 16'h1753; 14'h3112: x = 16'h1752; 14'h3113: x = 16'h1752; 14'h3114: x = 16'h1751; 14'h3115: x = 16'h1750; 14'h3116: x = 16'h174f; 14'h3117: x = 16'h174e; 14'h3118: x = 16'h174d; 14'h3119: x = 16'h174c; 14'h311a: x = 16'h174b; 14'h311b: x = 16'h174a; 14'h311c: x = 16'h1749; 14'h311d: x = 16'h1749; 14'h311e: x = 16'h1748; 14'h311f: x = 16'h1747; 14'h3120: x = 16'h1746; 14'h3121: x = 16'h1745; 14'h3122: x = 16'h1744; 14'h3123: x = 16'h1743; 14'h3124: x = 16'h1742; 14'h3125: x = 16'h1741; 14'h3126: x = 16'h1741; 14'h3127: x = 16'h1740; 14'h3128: x = 16'h173f; 14'h3129: x = 16'h173e; 14'h312a: x = 16'h173d; 14'h312b: x = 16'h173c; 14'h312c: x = 16'h173b; 14'h312d: x = 16'h173a; 14'h312e: x = 16'h1739; 14'h312f: x = 16'h1738; 14'h3130: x = 16'h1738; 14'h3131: x = 16'h1737; 14'h3132: x = 16'h1736; 14'h3133: x = 16'h1735; 14'h3134: x = 16'h1734; 14'h3135: x = 16'h1733; 14'h3136: x = 16'h1732; 14'h3137: x = 16'h1731; 14'h3138: x = 16'h1730; 14'h3139: x = 16'h172f; 14'h313a: x = 16'h172f; 14'h313b: x = 16'h172e; 14'h313c: x = 16'h172d; 14'h313d: x = 16'h172c; 14'h313e: x = 16'h172b; 14'h313f: x = 16'h172a; 14'h3140: x = 16'h1729; 14'h3141: x = 16'h1728; 14'h3142: x = 16'h1727; 14'h3143: x = 16'h1727; 14'h3144: x = 16'h1726; 14'h3145: x = 16'h1725; 14'h3146: x = 16'h1724; 14'h3147: x = 16'h1723; 14'h3148: x = 16'h1722; 14'h3149: x = 16'h1721; 14'h314a: x = 16'h1720; 14'h314b: x = 16'h171f; 14'h314c: x = 16'h171e; 14'h314d: x = 16'h171e; 14'h314e: x = 16'h171d; 14'h314f: x = 16'h171c; 14'h3150: x = 16'h171b; 14'h3151: x = 16'h171a; 14'h3152: x = 16'h1719; 14'h3153: x = 16'h1718; 14'h3154: x = 16'h1717; 14'h3155: x = 16'h1716; 14'h3156: x = 16'h1715; 14'h3157: x = 16'h1715; 14'h3158: x = 16'h1714; 14'h3159: x = 16'h1713; 14'h315a: x = 16'h1712; 14'h315b: x = 16'h1711; 14'h315c: x = 16'h1710; 14'h315d: x = 16'h170f; 14'h315e: x = 16'h170e; 14'h315f: x = 16'h170d; 14'h3160: x = 16'h170c; 14'h3161: x = 16'h170c; 14'h3162: x = 16'h170b; 14'h3163: x = 16'h170a; 14'h3164: x = 16'h1709; 14'h3165: x = 16'h1708; 14'h3166: x = 16'h1707; 14'h3167: x = 16'h1706; 14'h3168: x = 16'h1705; 14'h3169: x = 16'h1704; 14'h316a: x = 16'h1703; 14'h316b: x = 16'h1703; 14'h316c: x = 16'h1702; 14'h316d: x = 16'h1701; 14'h316e: x = 16'h1700; 14'h316f: x = 16'h16ff; 14'h3170: x = 16'h16fe; 14'h3171: x = 16'h16fd; 14'h3172: x = 16'h16fc; 14'h3173: x = 16'h16fb; 14'h3174: x = 16'h16fa; 14'h3175: x = 16'h16fa; 14'h3176: x = 16'h16f9; 14'h3177: x = 16'h16f8; 14'h3178: x = 16'h16f7; 14'h3179: x = 16'h16f6; 14'h317a: x = 16'h16f5; 14'h317b: x = 16'h16f4; 14'h317c: x = 16'h16f3; 14'h317d: x = 16'h16f2; 14'h317e: x = 16'h16f1; 14'h317f: x = 16'h16f1; 14'h3180: x = 16'h16f0; 14'h3181: x = 16'h16ef; 14'h3182: x = 16'h16ee; 14'h3183: x = 16'h16ed; 14'h3184: x = 16'h16ec; 14'h3185: x = 16'h16eb; 14'h3186: x = 16'h16ea; 14'h3187: x = 16'h16e9; 14'h3188: x = 16'h16e8; 14'h3189: x = 16'h16e8; 14'h318a: x = 16'h16e7; 14'h318b: x = 16'h16e6; 14'h318c: x = 16'h16e5; 14'h318d: x = 16'h16e4; 14'h318e: x = 16'h16e3; 14'h318f: x = 16'h16e2; 14'h3190: x = 16'h16e1; 14'h3191: x = 16'h16e0; 14'h3192: x = 16'h16df; 14'h3193: x = 16'h16de; 14'h3194: x = 16'h16de; 14'h3195: x = 16'h16dd; 14'h3196: x = 16'h16dc; 14'h3197: x = 16'h16db; 14'h3198: x = 16'h16da; 14'h3199: x = 16'h16d9; 14'h319a: x = 16'h16d8; 14'h319b: x = 16'h16d7; 14'h319c: x = 16'h16d6; 14'h319d: x = 16'h16d5; 14'h319e: x = 16'h16d5; 14'h319f: x = 16'h16d4; 14'h31a0: x = 16'h16d3; 14'h31a1: x = 16'h16d2; 14'h31a2: x = 16'h16d1; 14'h31a3: x = 16'h16d0; 14'h31a4: x = 16'h16cf; 14'h31a5: x = 16'h16ce; 14'h31a6: x = 16'h16cd; 14'h31a7: x = 16'h16cc; 14'h31a8: x = 16'h16cc; 14'h31a9: x = 16'h16cb; 14'h31aa: x = 16'h16ca; 14'h31ab: x = 16'h16c9; 14'h31ac: x = 16'h16c8; 14'h31ad: x = 16'h16c7; 14'h31ae: x = 16'h16c6; 14'h31af: x = 16'h16c5; 14'h31b0: x = 16'h16c4; 14'h31b1: x = 16'h16c3; 14'h31b2: x = 16'h16c2; 14'h31b3: x = 16'h16c2; 14'h31b4: x = 16'h16c1; 14'h31b5: x = 16'h16c0; 14'h31b6: x = 16'h16bf; 14'h31b7: x = 16'h16be; 14'h31b8: x = 16'h16bd; 14'h31b9: x = 16'h16bc; 14'h31ba: x = 16'h16bb; 14'h31bb: x = 16'h16ba; 14'h31bc: x = 16'h16b9; 14'h31bd: x = 16'h16b8; 14'h31be: x = 16'h16b8; 14'h31bf: x = 16'h16b7; 14'h31c0: x = 16'h16b6; 14'h31c1: x = 16'h16b5; 14'h31c2: x = 16'h16b4; 14'h31c3: x = 16'h16b3; 14'h31c4: x = 16'h16b2; 14'h31c5: x = 16'h16b1; 14'h31c6: x = 16'h16b0; 14'h31c7: x = 16'h16af; 14'h31c8: x = 16'h16af; 14'h31c9: x = 16'h16ae; 14'h31ca: x = 16'h16ad; 14'h31cb: x = 16'h16ac; 14'h31cc: x = 16'h16ab; 14'h31cd: x = 16'h16aa; 14'h31ce: x = 16'h16a9; 14'h31cf: x = 16'h16a8; 14'h31d0: x = 16'h16a7; 14'h31d1: x = 16'h16a6; 14'h31d2: x = 16'h16a5; 14'h31d3: x = 16'h16a5; 14'h31d4: x = 16'h16a4; 14'h31d5: x = 16'h16a3; 14'h31d6: x = 16'h16a2; 14'h31d7: x = 16'h16a1; 14'h31d8: x = 16'h16a0; 14'h31d9: x = 16'h169f; 14'h31da: x = 16'h169e; 14'h31db: x = 16'h169d; 14'h31dc: x = 16'h169c; 14'h31dd: x = 16'h169b; 14'h31de: x = 16'h169b; 14'h31df: x = 16'h169a; 14'h31e0: x = 16'h1699; 14'h31e1: x = 16'h1698; 14'h31e2: x = 16'h1697; 14'h31e3: x = 16'h1696; 14'h31e4: x = 16'h1695; 14'h31e5: x = 16'h1694; 14'h31e6: x = 16'h1693; 14'h31e7: x = 16'h1692; 14'h31e8: x = 16'h1691; 14'h31e9: x = 16'h1691; 14'h31ea: x = 16'h1690; 14'h31eb: x = 16'h168f; 14'h31ec: x = 16'h168e; 14'h31ed: x = 16'h168d; 14'h31ee: x = 16'h168c; 14'h31ef: x = 16'h168b; 14'h31f0: x = 16'h168a; 14'h31f1: x = 16'h1689; 14'h31f2: x = 16'h1688; 14'h31f3: x = 16'h1687; 14'h31f4: x = 16'h1687; 14'h31f5: x = 16'h1686; 14'h31f6: x = 16'h1685; 14'h31f7: x = 16'h1684; 14'h31f8: x = 16'h1683; 14'h31f9: x = 16'h1682; 14'h31fa: x = 16'h1681; 14'h31fb: x = 16'h1680; 14'h31fc: x = 16'h167f; 14'h31fd: x = 16'h167e; 14'h31fe: x = 16'h167d; 14'h31ff: x = 16'h167d; 14'h3200: x = 16'h167c; 14'h3201: x = 16'h167b; 14'h3202: x = 16'h167a; 14'h3203: x = 16'h1679; 14'h3204: x = 16'h1678; 14'h3205: x = 16'h1677; 14'h3206: x = 16'h1676; 14'h3207: x = 16'h1675; 14'h3208: x = 16'h1674; 14'h3209: x = 16'h1673; 14'h320a: x = 16'h1673; 14'h320b: x = 16'h1672; 14'h320c: x = 16'h1671; 14'h320d: x = 16'h1670; 14'h320e: x = 16'h166f; 14'h320f: x = 16'h166e; 14'h3210: x = 16'h166d; 14'h3211: x = 16'h166c; 14'h3212: x = 16'h166b; 14'h3213: x = 16'h166a; 14'h3214: x = 16'h1669; 14'h3215: x = 16'h1668; 14'h3216: x = 16'h1668; 14'h3217: x = 16'h1667; 14'h3218: x = 16'h1666; 14'h3219: x = 16'h1665; 14'h321a: x = 16'h1664; 14'h321b: x = 16'h1663; 14'h321c: x = 16'h1662; 14'h321d: x = 16'h1661; 14'h321e: x = 16'h1660; 14'h321f: x = 16'h165f; 14'h3220: x = 16'h165e; 14'h3221: x = 16'h165e; 14'h3222: x = 16'h165d; 14'h3223: x = 16'h165c; 14'h3224: x = 16'h165b; 14'h3225: x = 16'h165a; 14'h3226: x = 16'h1659; 14'h3227: x = 16'h1658; 14'h3228: x = 16'h1657; 14'h3229: x = 16'h1656; 14'h322a: x = 16'h1655; 14'h322b: x = 16'h1654; 14'h322c: x = 16'h1653; 14'h322d: x = 16'h1653; 14'h322e: x = 16'h1652; 14'h322f: x = 16'h1651; 14'h3230: x = 16'h1650; 14'h3231: x = 16'h164f; 14'h3232: x = 16'h164e; 14'h3233: x = 16'h164d; 14'h3234: x = 16'h164c; 14'h3235: x = 16'h164b; 14'h3236: x = 16'h164a; 14'h3237: x = 16'h1649; 14'h3238: x = 16'h1649; 14'h3239: x = 16'h1648; 14'h323a: x = 16'h1647; 14'h323b: x = 16'h1646; 14'h323c: x = 16'h1645; 14'h323d: x = 16'h1644; 14'h323e: x = 16'h1643; 14'h323f: x = 16'h1642; 14'h3240: x = 16'h1641; 14'h3241: x = 16'h1640; 14'h3242: x = 16'h163f; 14'h3243: x = 16'h163e; 14'h3244: x = 16'h163e; 14'h3245: x = 16'h163d; 14'h3246: x = 16'h163c; 14'h3247: x = 16'h163b; 14'h3248: x = 16'h163a; 14'h3249: x = 16'h1639; 14'h324a: x = 16'h1638; 14'h324b: x = 16'h1637; 14'h324c: x = 16'h1636; 14'h324d: x = 16'h1635; 14'h324e: x = 16'h1634; 14'h324f: x = 16'h1633; 14'h3250: x = 16'h1633; 14'h3251: x = 16'h1632; 14'h3252: x = 16'h1631; 14'h3253: x = 16'h1630; 14'h3254: x = 16'h162f; 14'h3255: x = 16'h162e; 14'h3256: x = 16'h162d; 14'h3257: x = 16'h162c; 14'h3258: x = 16'h162b; 14'h3259: x = 16'h162a; 14'h325a: x = 16'h1629; 14'h325b: x = 16'h1628; 14'h325c: x = 16'h1628; 14'h325d: x = 16'h1627; 14'h325e: x = 16'h1626; 14'h325f: x = 16'h1625; 14'h3260: x = 16'h1624; 14'h3261: x = 16'h1623; 14'h3262: x = 16'h1622; 14'h3263: x = 16'h1621; 14'h3264: x = 16'h1620; 14'h3265: x = 16'h161f; 14'h3266: x = 16'h161e; 14'h3267: x = 16'h161d; 14'h3268: x = 16'h161c; 14'h3269: x = 16'h161c; 14'h326a: x = 16'h161b; 14'h326b: x = 16'h161a; 14'h326c: x = 16'h1619; 14'h326d: x = 16'h1618; 14'h326e: x = 16'h1617; 14'h326f: x = 16'h1616; 14'h3270: x = 16'h1615; 14'h3271: x = 16'h1614; 14'h3272: x = 16'h1613; 14'h3273: x = 16'h1612; 14'h3274: x = 16'h1611; 14'h3275: x = 16'h1611; 14'h3276: x = 16'h1610; 14'h3277: x = 16'h160f; 14'h3278: x = 16'h160e; 14'h3279: x = 16'h160d; 14'h327a: x = 16'h160c; 14'h327b: x = 16'h160b; 14'h327c: x = 16'h160a; 14'h327d: x = 16'h1609; 14'h327e: x = 16'h1608; 14'h327f: x = 16'h1607; 14'h3280: x = 16'h1606; 14'h3281: x = 16'h1606; 14'h3282: x = 16'h1605; 14'h3283: x = 16'h1604; 14'h3284: x = 16'h1603; 14'h3285: x = 16'h1602; 14'h3286: x = 16'h1601; 14'h3287: x = 16'h1600; 14'h3288: x = 16'h15ff; 14'h3289: x = 16'h15fe; 14'h328a: x = 16'h15fd; 14'h328b: x = 16'h15fc; 14'h328c: x = 16'h15fb; 14'h328d: x = 16'h15fa; 14'h328e: x = 16'h15fa; 14'h328f: x = 16'h15f9; 14'h3290: x = 16'h15f8; 14'h3291: x = 16'h15f7; 14'h3292: x = 16'h15f6; 14'h3293: x = 16'h15f5; 14'h3294: x = 16'h15f4; 14'h3295: x = 16'h15f3; 14'h3296: x = 16'h15f2; 14'h3297: x = 16'h15f1; 14'h3298: x = 16'h15f0; 14'h3299: x = 16'h15ef; 14'h329a: x = 16'h15ee; 14'h329b: x = 16'h15ee; 14'h329c: x = 16'h15ed; 14'h329d: x = 16'h15ec; 14'h329e: x = 16'h15eb; 14'h329f: x = 16'h15ea; 14'h32a0: x = 16'h15e9; 14'h32a1: x = 16'h15e8; 14'h32a2: x = 16'h15e7; 14'h32a3: x = 16'h15e6; 14'h32a4: x = 16'h15e5; 14'h32a5: x = 16'h15e4; 14'h32a6: x = 16'h15e3; 14'h32a7: x = 16'h15e2; 14'h32a8: x = 16'h15e2; 14'h32a9: x = 16'h15e1; 14'h32aa: x = 16'h15e0; 14'h32ab: x = 16'h15df; 14'h32ac: x = 16'h15de; 14'h32ad: x = 16'h15dd; 14'h32ae: x = 16'h15dc; 14'h32af: x = 16'h15db; 14'h32b0: x = 16'h15da; 14'h32b1: x = 16'h15d9; 14'h32b2: x = 16'h15d8; 14'h32b3: x = 16'h15d7; 14'h32b4: x = 16'h15d6; 14'h32b5: x = 16'h15d6; 14'h32b6: x = 16'h15d5; 14'h32b7: x = 16'h15d4; 14'h32b8: x = 16'h15d3; 14'h32b9: x = 16'h15d2; 14'h32ba: x = 16'h15d1; 14'h32bb: x = 16'h15d0; 14'h32bc: x = 16'h15cf; 14'h32bd: x = 16'h15ce; 14'h32be: x = 16'h15cd; 14'h32bf: x = 16'h15cc; 14'h32c0: x = 16'h15cb; 14'h32c1: x = 16'h15ca; 14'h32c2: x = 16'h15c9; 14'h32c3: x = 16'h15c9; 14'h32c4: x = 16'h15c8; 14'h32c5: x = 16'h15c7; 14'h32c6: x = 16'h15c6; 14'h32c7: x = 16'h15c5; 14'h32c8: x = 16'h15c4; 14'h32c9: x = 16'h15c3; 14'h32ca: x = 16'h15c2; 14'h32cb: x = 16'h15c1; 14'h32cc: x = 16'h15c0; 14'h32cd: x = 16'h15bf; 14'h32ce: x = 16'h15be; 14'h32cf: x = 16'h15bd; 14'h32d0: x = 16'h15bd; 14'h32d1: x = 16'h15bc; 14'h32d2: x = 16'h15bb; 14'h32d3: x = 16'h15ba; 14'h32d4: x = 16'h15b9; 14'h32d5: x = 16'h15b8; 14'h32d6: x = 16'h15b7; 14'h32d7: x = 16'h15b6; 14'h32d8: x = 16'h15b5; 14'h32d9: x = 16'h15b4; 14'h32da: x = 16'h15b3; 14'h32db: x = 16'h15b2; 14'h32dc: x = 16'h15b1; 14'h32dd: x = 16'h15b0; 14'h32de: x = 16'h15b0; 14'h32df: x = 16'h15af; 14'h32e0: x = 16'h15ae; 14'h32e1: x = 16'h15ad; 14'h32e2: x = 16'h15ac; 14'h32e3: x = 16'h15ab; 14'h32e4: x = 16'h15aa; 14'h32e5: x = 16'h15a9; 14'h32e6: x = 16'h15a8; 14'h32e7: x = 16'h15a7; 14'h32e8: x = 16'h15a6; 14'h32e9: x = 16'h15a5; 14'h32ea: x = 16'h15a4; 14'h32eb: x = 16'h15a3; 14'h32ec: x = 16'h15a3; 14'h32ed: x = 16'h15a2; 14'h32ee: x = 16'h15a1; 14'h32ef: x = 16'h15a0; 14'h32f0: x = 16'h159f; 14'h32f1: x = 16'h159e; 14'h32f2: x = 16'h159d; 14'h32f3: x = 16'h159c; 14'h32f4: x = 16'h159b; 14'h32f5: x = 16'h159a; 14'h32f6: x = 16'h1599; 14'h32f7: x = 16'h1598; 14'h32f8: x = 16'h1597; 14'h32f9: x = 16'h1596; 14'h32fa: x = 16'h1596; 14'h32fb: x = 16'h1595; 14'h32fc: x = 16'h1594; 14'h32fd: x = 16'h1593; 14'h32fe: x = 16'h1592; 14'h32ff: x = 16'h1591; 14'h3300: x = 16'h1590; 14'h3301: x = 16'h158f; 14'h3302: x = 16'h158e; 14'h3303: x = 16'h158d; 14'h3304: x = 16'h158c; 14'h3305: x = 16'h158b; 14'h3306: x = 16'h158a; 14'h3307: x = 16'h1589; 14'h3308: x = 16'h1588; 14'h3309: x = 16'h1588; 14'h330a: x = 16'h1587; 14'h330b: x = 16'h1586; 14'h330c: x = 16'h1585; 14'h330d: x = 16'h1584; 14'h330e: x = 16'h1583; 14'h330f: x = 16'h1582; 14'h3310: x = 16'h1581; 14'h3311: x = 16'h1580; 14'h3312: x = 16'h157f; 14'h3313: x = 16'h157e; 14'h3314: x = 16'h157d; 14'h3315: x = 16'h157c; 14'h3316: x = 16'h157b; 14'h3317: x = 16'h157a; 14'h3318: x = 16'h157a; 14'h3319: x = 16'h1579; 14'h331a: x = 16'h1578; 14'h331b: x = 16'h1577; 14'h331c: x = 16'h1576; 14'h331d: x = 16'h1575; 14'h331e: x = 16'h1574; 14'h331f: x = 16'h1573; 14'h3320: x = 16'h1572; 14'h3321: x = 16'h1571; 14'h3322: x = 16'h1570; 14'h3323: x = 16'h156f; 14'h3324: x = 16'h156e; 14'h3325: x = 16'h156d; 14'h3326: x = 16'h156c; 14'h3327: x = 16'h156c; 14'h3328: x = 16'h156b; 14'h3329: x = 16'h156a; 14'h332a: x = 16'h1569; 14'h332b: x = 16'h1568; 14'h332c: x = 16'h1567; 14'h332d: x = 16'h1566; 14'h332e: x = 16'h1565; 14'h332f: x = 16'h1564; 14'h3330: x = 16'h1563; 14'h3331: x = 16'h1562; 14'h3332: x = 16'h1561; 14'h3333: x = 16'h1560; 14'h3334: x = 16'h155f; 14'h3335: x = 16'h155e; 14'h3336: x = 16'h155e; 14'h3337: x = 16'h155d; 14'h3338: x = 16'h155c; 14'h3339: x = 16'h155b; 14'h333a: x = 16'h155a; 14'h333b: x = 16'h1559; 14'h333c: x = 16'h1558; 14'h333d: x = 16'h1557; 14'h333e: x = 16'h1556; 14'h333f: x = 16'h1555; 14'h3340: x = 16'h1554; 14'h3341: x = 16'h1553; 14'h3342: x = 16'h1552; 14'h3343: x = 16'h1551; 14'h3344: x = 16'h1550; 14'h3345: x = 16'h154f; 14'h3346: x = 16'h154f; 14'h3347: x = 16'h154e; 14'h3348: x = 16'h154d; 14'h3349: x = 16'h154c; 14'h334a: x = 16'h154b; 14'h334b: x = 16'h154a; 14'h334c: x = 16'h1549; 14'h334d: x = 16'h1548; 14'h334e: x = 16'h1547; 14'h334f: x = 16'h1546; 14'h3350: x = 16'h1545; 14'h3351: x = 16'h1544; 14'h3352: x = 16'h1543; 14'h3353: x = 16'h1542; 14'h3354: x = 16'h1541; 14'h3355: x = 16'h1540; 14'h3356: x = 16'h1540; 14'h3357: x = 16'h153f; 14'h3358: x = 16'h153e; 14'h3359: x = 16'h153d; 14'h335a: x = 16'h153c; 14'h335b: x = 16'h153b; 14'h335c: x = 16'h153a; 14'h335d: x = 16'h1539; 14'h335e: x = 16'h1538; 14'h335f: x = 16'h1537; 14'h3360: x = 16'h1536; 14'h3361: x = 16'h1535; 14'h3362: x = 16'h1534; 14'h3363: x = 16'h1533; 14'h3364: x = 16'h1532; 14'h3365: x = 16'h1531; 14'h3366: x = 16'h1531; 14'h3367: x = 16'h1530; 14'h3368: x = 16'h152f; 14'h3369: x = 16'h152e; 14'h336a: x = 16'h152d; 14'h336b: x = 16'h152c; 14'h336c: x = 16'h152b; 14'h336d: x = 16'h152a; 14'h336e: x = 16'h1529; 14'h336f: x = 16'h1528; 14'h3370: x = 16'h1527; 14'h3371: x = 16'h1526; 14'h3372: x = 16'h1525; 14'h3373: x = 16'h1524; 14'h3374: x = 16'h1523; 14'h3375: x = 16'h1522; 14'h3376: x = 16'h1521; 14'h3377: x = 16'h1521; 14'h3378: x = 16'h1520; 14'h3379: x = 16'h151f; 14'h337a: x = 16'h151e; 14'h337b: x = 16'h151d; 14'h337c: x = 16'h151c; 14'h337d: x = 16'h151b; 14'h337e: x = 16'h151a; 14'h337f: x = 16'h1519; 14'h3380: x = 16'h1518; 14'h3381: x = 16'h1517; 14'h3382: x = 16'h1516; 14'h3383: x = 16'h1515; 14'h3384: x = 16'h1514; 14'h3385: x = 16'h1513; 14'h3386: x = 16'h1512; 14'h3387: x = 16'h1511; 14'h3388: x = 16'h1510; 14'h3389: x = 16'h1510; 14'h338a: x = 16'h150f; 14'h338b: x = 16'h150e; 14'h338c: x = 16'h150d; 14'h338d: x = 16'h150c; 14'h338e: x = 16'h150b; 14'h338f: x = 16'h150a; 14'h3390: x = 16'h1509; 14'h3391: x = 16'h1508; 14'h3392: x = 16'h1507; 14'h3393: x = 16'h1506; 14'h3394: x = 16'h1505; 14'h3395: x = 16'h1504; 14'h3396: x = 16'h1503; 14'h3397: x = 16'h1502; 14'h3398: x = 16'h1501; 14'h3399: x = 16'h1500; 14'h339a: x = 16'h14ff; 14'h339b: x = 16'h14ff; 14'h339c: x = 16'h14fe; 14'h339d: x = 16'h14fd; 14'h339e: x = 16'h14fc; 14'h339f: x = 16'h14fb; 14'h33a0: x = 16'h14fa; 14'h33a1: x = 16'h14f9; 14'h33a2: x = 16'h14f8; 14'h33a3: x = 16'h14f7; 14'h33a4: x = 16'h14f6; 14'h33a5: x = 16'h14f5; 14'h33a6: x = 16'h14f4; 14'h33a7: x = 16'h14f3; 14'h33a8: x = 16'h14f2; 14'h33a9: x = 16'h14f1; 14'h33aa: x = 16'h14f0; 14'h33ab: x = 16'h14ef; 14'h33ac: x = 16'h14ee; 14'h33ad: x = 16'h14ee; 14'h33ae: x = 16'h14ed; 14'h33af: x = 16'h14ec; 14'h33b0: x = 16'h14eb; 14'h33b1: x = 16'h14ea; 14'h33b2: x = 16'h14e9; 14'h33b3: x = 16'h14e8; 14'h33b4: x = 16'h14e7; 14'h33b5: x = 16'h14e6; 14'h33b6: x = 16'h14e5; 14'h33b7: x = 16'h14e4; 14'h33b8: x = 16'h14e3; 14'h33b9: x = 16'h14e2; 14'h33ba: x = 16'h14e1; 14'h33bb: x = 16'h14e0; 14'h33bc: x = 16'h14df; 14'h33bd: x = 16'h14de; 14'h33be: x = 16'h14dd; 14'h33bf: x = 16'h14dc; 14'h33c0: x = 16'h14dc; 14'h33c1: x = 16'h14db; 14'h33c2: x = 16'h14da; 14'h33c3: x = 16'h14d9; 14'h33c4: x = 16'h14d8; 14'h33c5: x = 16'h14d7; 14'h33c6: x = 16'h14d6; 14'h33c7: x = 16'h14d5; 14'h33c8: x = 16'h14d4; 14'h33c9: x = 16'h14d3; 14'h33ca: x = 16'h14d2; 14'h33cb: x = 16'h14d1; 14'h33cc: x = 16'h14d0; 14'h33cd: x = 16'h14cf; 14'h33ce: x = 16'h14ce; 14'h33cf: x = 16'h14cd; 14'h33d0: x = 16'h14cc; 14'h33d1: x = 16'h14cb; 14'h33d2: x = 16'h14ca; 14'h33d3: x = 16'h14c9; 14'h33d4: x = 16'h14c9; 14'h33d5: x = 16'h14c8; 14'h33d6: x = 16'h14c7; 14'h33d7: x = 16'h14c6; 14'h33d8: x = 16'h14c5; 14'h33d9: x = 16'h14c4; 14'h33da: x = 16'h14c3; 14'h33db: x = 16'h14c2; 14'h33dc: x = 16'h14c1; 14'h33dd: x = 16'h14c0; 14'h33de: x = 16'h14bf; 14'h33df: x = 16'h14be; 14'h33e0: x = 16'h14bd; 14'h33e1: x = 16'h14bc; 14'h33e2: x = 16'h14bb; 14'h33e3: x = 16'h14ba; 14'h33e4: x = 16'h14b9; 14'h33e5: x = 16'h14b8; 14'h33e6: x = 16'h14b7; 14'h33e7: x = 16'h14b6; 14'h33e8: x = 16'h14b5; 14'h33e9: x = 16'h14b5; 14'h33ea: x = 16'h14b4; 14'h33eb: x = 16'h14b3; 14'h33ec: x = 16'h14b2; 14'h33ed: x = 16'h14b1; 14'h33ee: x = 16'h14b0; 14'h33ef: x = 16'h14af; 14'h33f0: x = 16'h14ae; 14'h33f1: x = 16'h14ad; 14'h33f2: x = 16'h14ac; 14'h33f3: x = 16'h14ab; 14'h33f4: x = 16'h14aa; 14'h33f5: x = 16'h14a9; 14'h33f6: x = 16'h14a8; 14'h33f7: x = 16'h14a7; 14'h33f8: x = 16'h14a6; 14'h33f9: x = 16'h14a5; 14'h33fa: x = 16'h14a4; 14'h33fb: x = 16'h14a3; 14'h33fc: x = 16'h14a2; 14'h33fd: x = 16'h14a1; 14'h33fe: x = 16'h14a1; 14'h33ff: x = 16'h14a0; 14'h3400: x = 16'h149f; 14'h3401: x = 16'h149e; 14'h3402: x = 16'h149d; 14'h3403: x = 16'h149c; 14'h3404: x = 16'h149b; 14'h3405: x = 16'h149a; 14'h3406: x = 16'h1499; 14'h3407: x = 16'h1498; 14'h3408: x = 16'h1497; 14'h3409: x = 16'h1496; 14'h340a: x = 16'h1495; 14'h340b: x = 16'h1494; 14'h340c: x = 16'h1493; 14'h340d: x = 16'h1492; 14'h340e: x = 16'h1491; 14'h340f: x = 16'h1490; 14'h3410: x = 16'h148f; 14'h3411: x = 16'h148e; 14'h3412: x = 16'h148d; 14'h3413: x = 16'h148c; 14'h3414: x = 16'h148b; 14'h3415: x = 16'h148b; 14'h3416: x = 16'h148a; 14'h3417: x = 16'h1489; 14'h3418: x = 16'h1488; 14'h3419: x = 16'h1487; 14'h341a: x = 16'h1486; 14'h341b: x = 16'h1485; 14'h341c: x = 16'h1484; 14'h341d: x = 16'h1483; 14'h341e: x = 16'h1482; 14'h341f: x = 16'h1481; 14'h3420: x = 16'h1480; 14'h3421: x = 16'h147f; 14'h3422: x = 16'h147e; 14'h3423: x = 16'h147d; 14'h3424: x = 16'h147c; 14'h3425: x = 16'h147b; 14'h3426: x = 16'h147a; 14'h3427: x = 16'h1479; 14'h3428: x = 16'h1478; 14'h3429: x = 16'h1477; 14'h342a: x = 16'h1476; 14'h342b: x = 16'h1475; 14'h342c: x = 16'h1474; 14'h342d: x = 16'h1474; 14'h342e: x = 16'h1473; 14'h342f: x = 16'h1472; 14'h3430: x = 16'h1471; 14'h3431: x = 16'h1470; 14'h3432: x = 16'h146f; 14'h3433: x = 16'h146e; 14'h3434: x = 16'h146d; 14'h3435: x = 16'h146c; 14'h3436: x = 16'h146b; 14'h3437: x = 16'h146a; 14'h3438: x = 16'h1469; 14'h3439: x = 16'h1468; 14'h343a: x = 16'h1467; 14'h343b: x = 16'h1466; 14'h343c: x = 16'h1465; 14'h343d: x = 16'h1464; 14'h343e: x = 16'h1463; 14'h343f: x = 16'h1462; 14'h3440: x = 16'h1461; 14'h3441: x = 16'h1460; 14'h3442: x = 16'h145f; 14'h3443: x = 16'h145e; 14'h3444: x = 16'h145d; 14'h3445: x = 16'h145c; 14'h3446: x = 16'h145c; 14'h3447: x = 16'h145b; 14'h3448: x = 16'h145a; 14'h3449: x = 16'h1459; 14'h344a: x = 16'h1458; 14'h344b: x = 16'h1457; 14'h344c: x = 16'h1456; 14'h344d: x = 16'h1455; 14'h344e: x = 16'h1454; 14'h344f: x = 16'h1453; 14'h3450: x = 16'h1452; 14'h3451: x = 16'h1451; 14'h3452: x = 16'h1450; 14'h3453: x = 16'h144f; 14'h3454: x = 16'h144e; 14'h3455: x = 16'h144d; 14'h3456: x = 16'h144c; 14'h3457: x = 16'h144b; 14'h3458: x = 16'h144a; 14'h3459: x = 16'h1449; 14'h345a: x = 16'h1448; 14'h345b: x = 16'h1447; 14'h345c: x = 16'h1446; 14'h345d: x = 16'h1445; 14'h345e: x = 16'h1444; 14'h345f: x = 16'h1443; 14'h3460: x = 16'h1442; 14'h3461: x = 16'h1441; 14'h3462: x = 16'h1441; 14'h3463: x = 16'h1440; 14'h3464: x = 16'h143f; 14'h3465: x = 16'h143e; 14'h3466: x = 16'h143d; 14'h3467: x = 16'h143c; 14'h3468: x = 16'h143b; 14'h3469: x = 16'h143a; 14'h346a: x = 16'h1439; 14'h346b: x = 16'h1438; 14'h346c: x = 16'h1437; 14'h346d: x = 16'h1436; 14'h346e: x = 16'h1435; 14'h346f: x = 16'h1434; 14'h3470: x = 16'h1433; 14'h3471: x = 16'h1432; 14'h3472: x = 16'h1431; 14'h3473: x = 16'h1430; 14'h3474: x = 16'h142f; 14'h3475: x = 16'h142e; 14'h3476: x = 16'h142d; 14'h3477: x = 16'h142c; 14'h3478: x = 16'h142b; 14'h3479: x = 16'h142a; 14'h347a: x = 16'h1429; 14'h347b: x = 16'h1428; 14'h347c: x = 16'h1427; 14'h347d: x = 16'h1426; 14'h347e: x = 16'h1425; 14'h347f: x = 16'h1424; 14'h3480: x = 16'h1424; 14'h3481: x = 16'h1423; 14'h3482: x = 16'h1422; 14'h3483: x = 16'h1421; 14'h3484: x = 16'h1420; 14'h3485: x = 16'h141f; 14'h3486: x = 16'h141e; 14'h3487: x = 16'h141d; 14'h3488: x = 16'h141c; 14'h3489: x = 16'h141b; 14'h348a: x = 16'h141a; 14'h348b: x = 16'h1419; 14'h348c: x = 16'h1418; 14'h348d: x = 16'h1417; 14'h348e: x = 16'h1416; 14'h348f: x = 16'h1415; 14'h3490: x = 16'h1414; 14'h3491: x = 16'h1413; 14'h3492: x = 16'h1412; 14'h3493: x = 16'h1411; 14'h3494: x = 16'h1410; 14'h3495: x = 16'h140f; 14'h3496: x = 16'h140e; 14'h3497: x = 16'h140d; 14'h3498: x = 16'h140c; 14'h3499: x = 16'h140b; 14'h349a: x = 16'h140a; 14'h349b: x = 16'h1409; 14'h349c: x = 16'h1408; 14'h349d: x = 16'h1407; 14'h349e: x = 16'h1406; 14'h349f: x = 16'h1405; 14'h34a0: x = 16'h1404; 14'h34a1: x = 16'h1403; 14'h34a2: x = 16'h1403; 14'h34a3: x = 16'h1402; 14'h34a4: x = 16'h1401; 14'h34a5: x = 16'h1400; 14'h34a6: x = 16'h13ff; 14'h34a7: x = 16'h13fe; 14'h34a8: x = 16'h13fd; 14'h34a9: x = 16'h13fc; 14'h34aa: x = 16'h13fb; 14'h34ab: x = 16'h13fa; 14'h34ac: x = 16'h13f9; 14'h34ad: x = 16'h13f8; 14'h34ae: x = 16'h13f7; 14'h34af: x = 16'h13f6; 14'h34b0: x = 16'h13f5; 14'h34b1: x = 16'h13f4; 14'h34b2: x = 16'h13f3; 14'h34b3: x = 16'h13f2; 14'h34b4: x = 16'h13f1; 14'h34b5: x = 16'h13f0; 14'h34b6: x = 16'h13ef; 14'h34b7: x = 16'h13ee; 14'h34b8: x = 16'h13ed; 14'h34b9: x = 16'h13ec; 14'h34ba: x = 16'h13eb; 14'h34bb: x = 16'h13ea; 14'h34bc: x = 16'h13e9; 14'h34bd: x = 16'h13e8; 14'h34be: x = 16'h13e7; 14'h34bf: x = 16'h13e6; 14'h34c0: x = 16'h13e5; 14'h34c1: x = 16'h13e4; 14'h34c2: x = 16'h13e3; 14'h34c3: x = 16'h13e2; 14'h34c4: x = 16'h13e1; 14'h34c5: x = 16'h13e0; 14'h34c6: x = 16'h13df; 14'h34c7: x = 16'h13de; 14'h34c8: x = 16'h13dd; 14'h34c9: x = 16'h13dd; 14'h34ca: x = 16'h13dc; 14'h34cb: x = 16'h13db; 14'h34cc: x = 16'h13da; 14'h34cd: x = 16'h13d9; 14'h34ce: x = 16'h13d8; 14'h34cf: x = 16'h13d7; 14'h34d0: x = 16'h13d6; 14'h34d1: x = 16'h13d5; 14'h34d2: x = 16'h13d4; 14'h34d3: x = 16'h13d3; 14'h34d4: x = 16'h13d2; 14'h34d5: x = 16'h13d1; 14'h34d6: x = 16'h13d0; 14'h34d7: x = 16'h13cf; 14'h34d8: x = 16'h13ce; 14'h34d9: x = 16'h13cd; 14'h34da: x = 16'h13cc; 14'h34db: x = 16'h13cb; 14'h34dc: x = 16'h13ca; 14'h34dd: x = 16'h13c9; 14'h34de: x = 16'h13c8; 14'h34df: x = 16'h13c7; 14'h34e0: x = 16'h13c6; 14'h34e1: x = 16'h13c5; 14'h34e2: x = 16'h13c4; 14'h34e3: x = 16'h13c3; 14'h34e4: x = 16'h13c2; 14'h34e5: x = 16'h13c1; 14'h34e6: x = 16'h13c0; 14'h34e7: x = 16'h13bf; 14'h34e8: x = 16'h13be; 14'h34e9: x = 16'h13bd; 14'h34ea: x = 16'h13bc; 14'h34eb: x = 16'h13bb; 14'h34ec: x = 16'h13ba; 14'h34ed: x = 16'h13b9; 14'h34ee: x = 16'h13b8; 14'h34ef: x = 16'h13b7; 14'h34f0: x = 16'h13b6; 14'h34f1: x = 16'h13b5; 14'h34f2: x = 16'h13b4; 14'h34f3: x = 16'h13b3; 14'h34f4: x = 16'h13b2; 14'h34f5: x = 16'h13b1; 14'h34f6: x = 16'h13b0; 14'h34f7: x = 16'h13af; 14'h34f8: x = 16'h13ae; 14'h34f9: x = 16'h13ae; 14'h34fa: x = 16'h13ad; 14'h34fb: x = 16'h13ac; 14'h34fc: x = 16'h13ab; 14'h34fd: x = 16'h13aa; 14'h34fe: x = 16'h13a9; 14'h34ff: x = 16'h13a8; 14'h3500: x = 16'h13a7; 14'h3501: x = 16'h13a6; 14'h3502: x = 16'h13a5; 14'h3503: x = 16'h13a4; 14'h3504: x = 16'h13a3; 14'h3505: x = 16'h13a2; 14'h3506: x = 16'h13a1; 14'h3507: x = 16'h13a0; 14'h3508: x = 16'h139f; 14'h3509: x = 16'h139e; 14'h350a: x = 16'h139d; 14'h350b: x = 16'h139c; 14'h350c: x = 16'h139b; 14'h350d: x = 16'h139a; 14'h350e: x = 16'h1399; 14'h350f: x = 16'h1398; 14'h3510: x = 16'h1397; 14'h3511: x = 16'h1396; 14'h3512: x = 16'h1395; 14'h3513: x = 16'h1394; 14'h3514: x = 16'h1393; 14'h3515: x = 16'h1392; 14'h3516: x = 16'h1391; 14'h3517: x = 16'h1390; 14'h3518: x = 16'h138f; 14'h3519: x = 16'h138e; 14'h351a: x = 16'h138d; 14'h351b: x = 16'h138c; 14'h351c: x = 16'h138b; 14'h351d: x = 16'h138a; 14'h351e: x = 16'h1389; 14'h351f: x = 16'h1388; 14'h3520: x = 16'h1387; 14'h3521: x = 16'h1386; 14'h3522: x = 16'h1385; 14'h3523: x = 16'h1384; 14'h3524: x = 16'h1383; 14'h3525: x = 16'h1382; 14'h3526: x = 16'h1381; 14'h3527: x = 16'h1380; 14'h3528: x = 16'h137f; 14'h3529: x = 16'h137e; 14'h352a: x = 16'h137d; 14'h352b: x = 16'h137c; 14'h352c: x = 16'h137b; 14'h352d: x = 16'h137a; 14'h352e: x = 16'h1379; 14'h352f: x = 16'h1378; 14'h3530: x = 16'h1377; 14'h3531: x = 16'h1376; 14'h3532: x = 16'h1375; 14'h3533: x = 16'h1374; 14'h3534: x = 16'h1373; 14'h3535: x = 16'h1372; 14'h3536: x = 16'h1371; 14'h3537: x = 16'h1370; 14'h3538: x = 16'h136f; 14'h3539: x = 16'h136e; 14'h353a: x = 16'h136d; 14'h353b: x = 16'h136c; 14'h353c: x = 16'h136b; 14'h353d: x = 16'h136a; 14'h353e: x = 16'h1369; 14'h353f: x = 16'h1368; 14'h3540: x = 16'h1367; 14'h3541: x = 16'h1366; 14'h3542: x = 16'h1365; 14'h3543: x = 16'h1364; 14'h3544: x = 16'h1363; 14'h3545: x = 16'h1363; 14'h3546: x = 16'h1362; 14'h3547: x = 16'h1361; 14'h3548: x = 16'h1360; 14'h3549: x = 16'h135f; 14'h354a: x = 16'h135e; 14'h354b: x = 16'h135d; 14'h354c: x = 16'h135c; 14'h354d: x = 16'h135b; 14'h354e: x = 16'h135a; 14'h354f: x = 16'h1359; 14'h3550: x = 16'h1358; 14'h3551: x = 16'h1357; 14'h3552: x = 16'h1356; 14'h3553: x = 16'h1355; 14'h3554: x = 16'h1354; 14'h3555: x = 16'h1353; 14'h3556: x = 16'h1352; 14'h3557: x = 16'h1351; 14'h3558: x = 16'h1350; 14'h3559: x = 16'h134f; 14'h355a: x = 16'h134e; 14'h355b: x = 16'h134d; 14'h355c: x = 16'h134c; 14'h355d: x = 16'h134b; 14'h355e: x = 16'h134a; 14'h355f: x = 16'h1349; 14'h3560: x = 16'h1348; 14'h3561: x = 16'h1347; 14'h3562: x = 16'h1346; 14'h3563: x = 16'h1345; 14'h3564: x = 16'h1344; 14'h3565: x = 16'h1343; 14'h3566: x = 16'h1342; 14'h3567: x = 16'h1341; 14'h3568: x = 16'h1340; 14'h3569: x = 16'h133f; 14'h356a: x = 16'h133e; 14'h356b: x = 16'h133d; 14'h356c: x = 16'h133c; 14'h356d: x = 16'h133b; 14'h356e: x = 16'h133a; 14'h356f: x = 16'h1339; 14'h3570: x = 16'h1338; 14'h3571: x = 16'h1337; 14'h3572: x = 16'h1336; 14'h3573: x = 16'h1335; 14'h3574: x = 16'h1334; 14'h3575: x = 16'h1333; 14'h3576: x = 16'h1332; 14'h3577: x = 16'h1331; 14'h3578: x = 16'h1330; 14'h3579: x = 16'h132f; 14'h357a: x = 16'h132e; 14'h357b: x = 16'h132d; 14'h357c: x = 16'h132c; 14'h357d: x = 16'h132b; 14'h357e: x = 16'h132a; 14'h357f: x = 16'h1329; 14'h3580: x = 16'h1328; 14'h3581: x = 16'h1327; 14'h3582: x = 16'h1326; 14'h3583: x = 16'h1325; 14'h3584: x = 16'h1324; 14'h3585: x = 16'h1323; 14'h3586: x = 16'h1322; 14'h3587: x = 16'h1321; 14'h3588: x = 16'h1320; 14'h3589: x = 16'h131f; 14'h358a: x = 16'h131e; 14'h358b: x = 16'h131d; 14'h358c: x = 16'h131c; 14'h358d: x = 16'h131b; 14'h358e: x = 16'h131a; 14'h358f: x = 16'h1319; 14'h3590: x = 16'h1318; 14'h3591: x = 16'h1317; 14'h3592: x = 16'h1316; 14'h3593: x = 16'h1315; 14'h3594: x = 16'h1314; 14'h3595: x = 16'h1313; 14'h3596: x = 16'h1312; 14'h3597: x = 16'h1311; 14'h3598: x = 16'h1310; 14'h3599: x = 16'h130f; 14'h359a: x = 16'h130e; 14'h359b: x = 16'h130d; 14'h359c: x = 16'h130c; 14'h359d: x = 16'h130b; 14'h359e: x = 16'h130a; 14'h359f: x = 16'h1309; 14'h35a0: x = 16'h1308; 14'h35a1: x = 16'h1307; 14'h35a2: x = 16'h1306; 14'h35a3: x = 16'h1305; 14'h35a4: x = 16'h1304; 14'h35a5: x = 16'h1303; 14'h35a6: x = 16'h1302; 14'h35a7: x = 16'h1301; 14'h35a8: x = 16'h1300; 14'h35a9: x = 16'h12ff; 14'h35aa: x = 16'h12fe; 14'h35ab: x = 16'h12fd; 14'h35ac: x = 16'h12fc; 14'h35ad: x = 16'h12fb; 14'h35ae: x = 16'h12fa; 14'h35af: x = 16'h12f9; 14'h35b0: x = 16'h12f8; 14'h35b1: x = 16'h12f7; 14'h35b2: x = 16'h12f6; 14'h35b3: x = 16'h12f5; 14'h35b4: x = 16'h12f4; 14'h35b5: x = 16'h12f3; 14'h35b6: x = 16'h12f2; 14'h35b7: x = 16'h12f1; 14'h35b8: x = 16'h12f0; 14'h35b9: x = 16'h12ef; 14'h35ba: x = 16'h12ee; 14'h35bb: x = 16'h12ed; 14'h35bc: x = 16'h12ec; 14'h35bd: x = 16'h12eb; 14'h35be: x = 16'h12ea; 14'h35bf: x = 16'h12e9; 14'h35c0: x = 16'h12e8; 14'h35c1: x = 16'h12e7; 14'h35c2: x = 16'h12e6; 14'h35c3: x = 16'h12e5; 14'h35c4: x = 16'h12e4; 14'h35c5: x = 16'h12e3; 14'h35c6: x = 16'h12e2; 14'h35c7: x = 16'h12e1; 14'h35c8: x = 16'h12e0; 14'h35c9: x = 16'h12de; 14'h35ca: x = 16'h12dd; 14'h35cb: x = 16'h12dc; 14'h35cc: x = 16'h12db; 14'h35cd: x = 16'h12da; 14'h35ce: x = 16'h12d9; 14'h35cf: x = 16'h12d8; 14'h35d0: x = 16'h12d7; 14'h35d1: x = 16'h12d6; 14'h35d2: x = 16'h12d5; 14'h35d3: x = 16'h12d4; 14'h35d4: x = 16'h12d3; 14'h35d5: x = 16'h12d2; 14'h35d6: x = 16'h12d1; 14'h35d7: x = 16'h12d0; 14'h35d8: x = 16'h12cf; 14'h35d9: x = 16'h12ce; 14'h35da: x = 16'h12cd; 14'h35db: x = 16'h12cc; 14'h35dc: x = 16'h12cb; 14'h35dd: x = 16'h12ca; 14'h35de: x = 16'h12c9; 14'h35df: x = 16'h12c8; 14'h35e0: x = 16'h12c7; 14'h35e1: x = 16'h12c6; 14'h35e2: x = 16'h12c5; 14'h35e3: x = 16'h12c4; 14'h35e4: x = 16'h12c3; 14'h35e5: x = 16'h12c2; 14'h35e6: x = 16'h12c1; 14'h35e7: x = 16'h12c0; 14'h35e8: x = 16'h12bf; 14'h35e9: x = 16'h12be; 14'h35ea: x = 16'h12bd; 14'h35eb: x = 16'h12bc; 14'h35ec: x = 16'h12bb; 14'h35ed: x = 16'h12ba; 14'h35ee: x = 16'h12b9; 14'h35ef: x = 16'h12b8; 14'h35f0: x = 16'h12b7; 14'h35f1: x = 16'h12b6; 14'h35f2: x = 16'h12b5; 14'h35f3: x = 16'h12b4; 14'h35f4: x = 16'h12b3; 14'h35f5: x = 16'h12b2; 14'h35f6: x = 16'h12b1; 14'h35f7: x = 16'h12b0; 14'h35f8: x = 16'h12af; 14'h35f9: x = 16'h12ae; 14'h35fa: x = 16'h12ad; 14'h35fb: x = 16'h12ac; 14'h35fc: x = 16'h12ab; 14'h35fd: x = 16'h12aa; 14'h35fe: x = 16'h12a9; 14'h35ff: x = 16'h12a8; 14'h3600: x = 16'h12a7; 14'h3601: x = 16'h12a6; 14'h3602: x = 16'h12a5; 14'h3603: x = 16'h12a4; 14'h3604: x = 16'h12a3; 14'h3605: x = 16'h12a2; 14'h3606: x = 16'h12a1; 14'h3607: x = 16'h12a0; 14'h3608: x = 16'h129f; 14'h3609: x = 16'h129e; 14'h360a: x = 16'h129d; 14'h360b: x = 16'h129c; 14'h360c: x = 16'h129b; 14'h360d: x = 16'h129a; 14'h360e: x = 16'h1299; 14'h360f: x = 16'h1298; 14'h3610: x = 16'h1297; 14'h3611: x = 16'h1295; 14'h3612: x = 16'h1294; 14'h3613: x = 16'h1293; 14'h3614: x = 16'h1292; 14'h3615: x = 16'h1291; 14'h3616: x = 16'h1290; 14'h3617: x = 16'h128f; 14'h3618: x = 16'h128e; 14'h3619: x = 16'h128d; 14'h361a: x = 16'h128c; 14'h361b: x = 16'h128b; 14'h361c: x = 16'h128a; 14'h361d: x = 16'h1289; 14'h361e: x = 16'h1288; 14'h361f: x = 16'h1287; 14'h3620: x = 16'h1286; 14'h3621: x = 16'h1285; 14'h3622: x = 16'h1284; 14'h3623: x = 16'h1283; 14'h3624: x = 16'h1282; 14'h3625: x = 16'h1281; 14'h3626: x = 16'h1280; 14'h3627: x = 16'h127f; 14'h3628: x = 16'h127e; 14'h3629: x = 16'h127d; 14'h362a: x = 16'h127c; 14'h362b: x = 16'h127b; 14'h362c: x = 16'h127a; 14'h362d: x = 16'h1279; 14'h362e: x = 16'h1278; 14'h362f: x = 16'h1277; 14'h3630: x = 16'h1276; 14'h3631: x = 16'h1275; 14'h3632: x = 16'h1274; 14'h3633: x = 16'h1273; 14'h3634: x = 16'h1272; 14'h3635: x = 16'h1271; 14'h3636: x = 16'h1270; 14'h3637: x = 16'h126f; 14'h3638: x = 16'h126e; 14'h3639: x = 16'h126d; 14'h363a: x = 16'h126c; 14'h363b: x = 16'h126b; 14'h363c: x = 16'h126a; 14'h363d: x = 16'h1269; 14'h363e: x = 16'h1267; 14'h363f: x = 16'h1266; 14'h3640: x = 16'h1265; 14'h3641: x = 16'h1264; 14'h3642: x = 16'h1263; 14'h3643: x = 16'h1262; 14'h3644: x = 16'h1261; 14'h3645: x = 16'h1260; 14'h3646: x = 16'h125f; 14'h3647: x = 16'h125e; 14'h3648: x = 16'h125d; 14'h3649: x = 16'h125c; 14'h364a: x = 16'h125b; 14'h364b: x = 16'h125a; 14'h364c: x = 16'h1259; 14'h364d: x = 16'h1258; 14'h364e: x = 16'h1257; 14'h364f: x = 16'h1256; 14'h3650: x = 16'h1255; 14'h3651: x = 16'h1254; 14'h3652: x = 16'h1253; 14'h3653: x = 16'h1252; 14'h3654: x = 16'h1251; 14'h3655: x = 16'h1250; 14'h3656: x = 16'h124f; 14'h3657: x = 16'h124e; 14'h3658: x = 16'h124d; 14'h3659: x = 16'h124c; 14'h365a: x = 16'h124b; 14'h365b: x = 16'h124a; 14'h365c: x = 16'h1249; 14'h365d: x = 16'h1248; 14'h365e: x = 16'h1247; 14'h365f: x = 16'h1246; 14'h3660: x = 16'h1245; 14'h3661: x = 16'h1243; 14'h3662: x = 16'h1242; 14'h3663: x = 16'h1241; 14'h3664: x = 16'h1240; 14'h3665: x = 16'h123f; 14'h3666: x = 16'h123e; 14'h3667: x = 16'h123d; 14'h3668: x = 16'h123c; 14'h3669: x = 16'h123b; 14'h366a: x = 16'h123a; 14'h366b: x = 16'h1239; 14'h366c: x = 16'h1238; 14'h366d: x = 16'h1237; 14'h366e: x = 16'h1236; 14'h366f: x = 16'h1235; 14'h3670: x = 16'h1234; 14'h3671: x = 16'h1233; 14'h3672: x = 16'h1232; 14'h3673: x = 16'h1231; 14'h3674: x = 16'h1230; 14'h3675: x = 16'h122f; 14'h3676: x = 16'h122e; 14'h3677: x = 16'h122d; 14'h3678: x = 16'h122c; 14'h3679: x = 16'h122b; 14'h367a: x = 16'h122a; 14'h367b: x = 16'h1229; 14'h367c: x = 16'h1228; 14'h367d: x = 16'h1227; 14'h367e: x = 16'h1226; 14'h367f: x = 16'h1225; 14'h3680: x = 16'h1223; 14'h3681: x = 16'h1222; 14'h3682: x = 16'h1221; 14'h3683: x = 16'h1220; 14'h3684: x = 16'h121f; 14'h3685: x = 16'h121e; 14'h3686: x = 16'h121d; 14'h3687: x = 16'h121c; 14'h3688: x = 16'h121b; 14'h3689: x = 16'h121a; 14'h368a: x = 16'h1219; 14'h368b: x = 16'h1218; 14'h368c: x = 16'h1217; 14'h368d: x = 16'h1216; 14'h368e: x = 16'h1215; 14'h368f: x = 16'h1214; 14'h3690: x = 16'h1213; 14'h3691: x = 16'h1212; 14'h3692: x = 16'h1211; 14'h3693: x = 16'h1210; 14'h3694: x = 16'h120f; 14'h3695: x = 16'h120e; 14'h3696: x = 16'h120d; 14'h3697: x = 16'h120c; 14'h3698: x = 16'h120b; 14'h3699: x = 16'h120a; 14'h369a: x = 16'h1208; 14'h369b: x = 16'h1207; 14'h369c: x = 16'h1206; 14'h369d: x = 16'h1205; 14'h369e: x = 16'h1204; 14'h369f: x = 16'h1203; 14'h36a0: x = 16'h1202; 14'h36a1: x = 16'h1201; 14'h36a2: x = 16'h1200; 14'h36a3: x = 16'h11ff; 14'h36a4: x = 16'h11fe; 14'h36a5: x = 16'h11fd; 14'h36a6: x = 16'h11fc; 14'h36a7: x = 16'h11fb; 14'h36a8: x = 16'h11fa; 14'h36a9: x = 16'h11f9; 14'h36aa: x = 16'h11f8; 14'h36ab: x = 16'h11f7; 14'h36ac: x = 16'h11f6; 14'h36ad: x = 16'h11f5; 14'h36ae: x = 16'h11f4; 14'h36af: x = 16'h11f3; 14'h36b0: x = 16'h11f2; 14'h36b1: x = 16'h11f1; 14'h36b2: x = 16'h11ef; 14'h36b3: x = 16'h11ee; 14'h36b4: x = 16'h11ed; 14'h36b5: x = 16'h11ec; 14'h36b6: x = 16'h11eb; 14'h36b7: x = 16'h11ea; 14'h36b8: x = 16'h11e9; 14'h36b9: x = 16'h11e8; 14'h36ba: x = 16'h11e7; 14'h36bb: x = 16'h11e6; 14'h36bc: x = 16'h11e5; 14'h36bd: x = 16'h11e4; 14'h36be: x = 16'h11e3; 14'h36bf: x = 16'h11e2; 14'h36c0: x = 16'h11e1; 14'h36c1: x = 16'h11e0; 14'h36c2: x = 16'h11df; 14'h36c3: x = 16'h11de; 14'h36c4: x = 16'h11dd; 14'h36c5: x = 16'h11dc; 14'h36c6: x = 16'h11db; 14'h36c7: x = 16'h11da; 14'h36c8: x = 16'h11d8; 14'h36c9: x = 16'h11d7; 14'h36ca: x = 16'h11d6; 14'h36cb: x = 16'h11d5; 14'h36cc: x = 16'h11d4; 14'h36cd: x = 16'h11d3; 14'h36ce: x = 16'h11d2; 14'h36cf: x = 16'h11d1; 14'h36d0: x = 16'h11d0; 14'h36d1: x = 16'h11cf; 14'h36d2: x = 16'h11ce; 14'h36d3: x = 16'h11cd; 14'h36d4: x = 16'h11cc; 14'h36d5: x = 16'h11cb; 14'h36d6: x = 16'h11ca; 14'h36d7: x = 16'h11c9; 14'h36d8: x = 16'h11c8; 14'h36d9: x = 16'h11c7; 14'h36da: x = 16'h11c6; 14'h36db: x = 16'h11c5; 14'h36dc: x = 16'h11c3; 14'h36dd: x = 16'h11c2; 14'h36de: x = 16'h11c1; 14'h36df: x = 16'h11c0; 14'h36e0: x = 16'h11bf; 14'h36e1: x = 16'h11be; 14'h36e2: x = 16'h11bd; 14'h36e3: x = 16'h11bc; 14'h36e4: x = 16'h11bb; 14'h36e5: x = 16'h11ba; 14'h36e6: x = 16'h11b9; 14'h36e7: x = 16'h11b8; 14'h36e8: x = 16'h11b7; 14'h36e9: x = 16'h11b6; 14'h36ea: x = 16'h11b5; 14'h36eb: x = 16'h11b4; 14'h36ec: x = 16'h11b3; 14'h36ed: x = 16'h11b2; 14'h36ee: x = 16'h11b1; 14'h36ef: x = 16'h11b0; 14'h36f0: x = 16'h11ae; 14'h36f1: x = 16'h11ad; 14'h36f2: x = 16'h11ac; 14'h36f3: x = 16'h11ab; 14'h36f4: x = 16'h11aa; 14'h36f5: x = 16'h11a9; 14'h36f6: x = 16'h11a8; 14'h36f7: x = 16'h11a7; 14'h36f8: x = 16'h11a6; 14'h36f9: x = 16'h11a5; 14'h36fa: x = 16'h11a4; 14'h36fb: x = 16'h11a3; 14'h36fc: x = 16'h11a2; 14'h36fd: x = 16'h11a1; 14'h36fe: x = 16'h11a0; 14'h36ff: x = 16'h119f; 14'h3700: x = 16'h119e; 14'h3701: x = 16'h119d; 14'h3702: x = 16'h119b; 14'h3703: x = 16'h119a; 14'h3704: x = 16'h1199; 14'h3705: x = 16'h1198; 14'h3706: x = 16'h1197; 14'h3707: x = 16'h1196; 14'h3708: x = 16'h1195; 14'h3709: x = 16'h1194; 14'h370a: x = 16'h1193; 14'h370b: x = 16'h1192; 14'h370c: x = 16'h1191; 14'h370d: x = 16'h1190; 14'h370e: x = 16'h118f; 14'h370f: x = 16'h118e; 14'h3710: x = 16'h118d; 14'h3711: x = 16'h118c; 14'h3712: x = 16'h118b; 14'h3713: x = 16'h1189; 14'h3714: x = 16'h1188; 14'h3715: x = 16'h1187; 14'h3716: x = 16'h1186; 14'h3717: x = 16'h1185; 14'h3718: x = 16'h1184; 14'h3719: x = 16'h1183; 14'h371a: x = 16'h1182; 14'h371b: x = 16'h1181; 14'h371c: x = 16'h1180; 14'h371d: x = 16'h117f; 14'h371e: x = 16'h117e; 14'h371f: x = 16'h117d; 14'h3720: x = 16'h117c; 14'h3721: x = 16'h117b; 14'h3722: x = 16'h117a; 14'h3723: x = 16'h1178; 14'h3724: x = 16'h1177; 14'h3725: x = 16'h1176; 14'h3726: x = 16'h1175; 14'h3727: x = 16'h1174; 14'h3728: x = 16'h1173; 14'h3729: x = 16'h1172; 14'h372a: x = 16'h1171; 14'h372b: x = 16'h1170; 14'h372c: x = 16'h116f; 14'h372d: x = 16'h116e; 14'h372e: x = 16'h116d; 14'h372f: x = 16'h116c; 14'h3730: x = 16'h116b; 14'h3731: x = 16'h116a; 14'h3732: x = 16'h1169; 14'h3733: x = 16'h1167; 14'h3734: x = 16'h1166; 14'h3735: x = 16'h1165; 14'h3736: x = 16'h1164; 14'h3737: x = 16'h1163; 14'h3738: x = 16'h1162; 14'h3739: x = 16'h1161; 14'h373a: x = 16'h1160; 14'h373b: x = 16'h115f; 14'h373c: x = 16'h115e; 14'h373d: x = 16'h115d; 14'h373e: x = 16'h115c; 14'h373f: x = 16'h115b; 14'h3740: x = 16'h115a; 14'h3741: x = 16'h1159; 14'h3742: x = 16'h1157; 14'h3743: x = 16'h1156; 14'h3744: x = 16'h1155; 14'h3745: x = 16'h1154; 14'h3746: x = 16'h1153; 14'h3747: x = 16'h1152; 14'h3748: x = 16'h1151; 14'h3749: x = 16'h1150; 14'h374a: x = 16'h114f; 14'h374b: x = 16'h114e; 14'h374c: x = 16'h114d; 14'h374d: x = 16'h114c; 14'h374e: x = 16'h114b; 14'h374f: x = 16'h114a; 14'h3750: x = 16'h1148; 14'h3751: x = 16'h1147; 14'h3752: x = 16'h1146; 14'h3753: x = 16'h1145; 14'h3754: x = 16'h1144; 14'h3755: x = 16'h1143; 14'h3756: x = 16'h1142; 14'h3757: x = 16'h1141; 14'h3758: x = 16'h1140; 14'h3759: x = 16'h113f; 14'h375a: x = 16'h113e; 14'h375b: x = 16'h113d; 14'h375c: x = 16'h113c; 14'h375d: x = 16'h113b; 14'h375e: x = 16'h1139; 14'h375f: x = 16'h1138; 14'h3760: x = 16'h1137; 14'h3761: x = 16'h1136; 14'h3762: x = 16'h1135; 14'h3763: x = 16'h1134; 14'h3764: x = 16'h1133; 14'h3765: x = 16'h1132; 14'h3766: x = 16'h1131; 14'h3767: x = 16'h1130; 14'h3768: x = 16'h112f; 14'h3769: x = 16'h112e; 14'h376a: x = 16'h112d; 14'h376b: x = 16'h112b; 14'h376c: x = 16'h112a; 14'h376d: x = 16'h1129; 14'h376e: x = 16'h1128; 14'h376f: x = 16'h1127; 14'h3770: x = 16'h1126; 14'h3771: x = 16'h1125; 14'h3772: x = 16'h1124; 14'h3773: x = 16'h1123; 14'h3774: x = 16'h1122; 14'h3775: x = 16'h1121; 14'h3776: x = 16'h1120; 14'h3777: x = 16'h111f; 14'h3778: x = 16'h111d; 14'h3779: x = 16'h111c; 14'h377a: x = 16'h111b; 14'h377b: x = 16'h111a; 14'h377c: x = 16'h1119; 14'h377d: x = 16'h1118; 14'h377e: x = 16'h1117; 14'h377f: x = 16'h1116; 14'h3780: x = 16'h1115; 14'h3781: x = 16'h1114; 14'h3782: x = 16'h1113; 14'h3783: x = 16'h1112; 14'h3784: x = 16'h1111; 14'h3785: x = 16'h110f; 14'h3786: x = 16'h110e; 14'h3787: x = 16'h110d; 14'h3788: x = 16'h110c; 14'h3789: x = 16'h110b; 14'h378a: x = 16'h110a; 14'h378b: x = 16'h1109; 14'h378c: x = 16'h1108; 14'h378d: x = 16'h1107; 14'h378e: x = 16'h1106; 14'h378f: x = 16'h1105; 14'h3790: x = 16'h1104; 14'h3791: x = 16'h1102; 14'h3792: x = 16'h1101; 14'h3793: x = 16'h1100; 14'h3794: x = 16'h10ff; 14'h3795: x = 16'h10fe; 14'h3796: x = 16'h10fd; 14'h3797: x = 16'h10fc; 14'h3798: x = 16'h10fb; 14'h3799: x = 16'h10fa; 14'h379a: x = 16'h10f9; 14'h379b: x = 16'h10f8; 14'h379c: x = 16'h10f7; 14'h379d: x = 16'h10f5; 14'h379e: x = 16'h10f4; 14'h379f: x = 16'h10f3; 14'h37a0: x = 16'h10f2; 14'h37a1: x = 16'h10f1; 14'h37a2: x = 16'h10f0; 14'h37a3: x = 16'h10ef; 14'h37a4: x = 16'h10ee; 14'h37a5: x = 16'h10ed; 14'h37a6: x = 16'h10ec; 14'h37a7: x = 16'h10eb; 14'h37a8: x = 16'h10e9; 14'h37a9: x = 16'h10e8; 14'h37aa: x = 16'h10e7; 14'h37ab: x = 16'h10e6; 14'h37ac: x = 16'h10e5; 14'h37ad: x = 16'h10e4; 14'h37ae: x = 16'h10e3; 14'h37af: x = 16'h10e2; 14'h37b0: x = 16'h10e1; 14'h37b1: x = 16'h10e0; 14'h37b2: x = 16'h10df; 14'h37b3: x = 16'h10dd; 14'h37b4: x = 16'h10dc; 14'h37b5: x = 16'h10db; 14'h37b6: x = 16'h10da; 14'h37b7: x = 16'h10d9; 14'h37b8: x = 16'h10d8; 14'h37b9: x = 16'h10d7; 14'h37ba: x = 16'h10d6; 14'h37bb: x = 16'h10d5; 14'h37bc: x = 16'h10d4; 14'h37bd: x = 16'h10d3; 14'h37be: x = 16'h10d1; 14'h37bf: x = 16'h10d0; 14'h37c0: x = 16'h10cf; 14'h37c1: x = 16'h10ce; 14'h37c2: x = 16'h10cd; 14'h37c3: x = 16'h10cc; 14'h37c4: x = 16'h10cb; 14'h37c5: x = 16'h10ca; 14'h37c6: x = 16'h10c9; 14'h37c7: x = 16'h10c8; 14'h37c8: x = 16'h10c7; 14'h37c9: x = 16'h10c5; 14'h37ca: x = 16'h10c4; 14'h37cb: x = 16'h10c3; 14'h37cc: x = 16'h10c2; 14'h37cd: x = 16'h10c1; 14'h37ce: x = 16'h10c0; 14'h37cf: x = 16'h10bf; 14'h37d0: x = 16'h10be; 14'h37d1: x = 16'h10bd; 14'h37d2: x = 16'h10bc; 14'h37d3: x = 16'h10bb; 14'h37d4: x = 16'h10b9; 14'h37d5: x = 16'h10b8; 14'h37d6: x = 16'h10b7; 14'h37d7: x = 16'h10b6; 14'h37d8: x = 16'h10b5; 14'h37d9: x = 16'h10b4; 14'h37da: x = 16'h10b3; 14'h37db: x = 16'h10b2; 14'h37dc: x = 16'h10b1; 14'h37dd: x = 16'h10b0; 14'h37de: x = 16'h10ae; 14'h37df: x = 16'h10ad; 14'h37e0: x = 16'h10ac; 14'h37e1: x = 16'h10ab; 14'h37e2: x = 16'h10aa; 14'h37e3: x = 16'h10a9; 14'h37e4: x = 16'h10a8; 14'h37e5: x = 16'h10a7; 14'h37e6: x = 16'h10a6; 14'h37e7: x = 16'h10a5; 14'h37e8: x = 16'h10a3; 14'h37e9: x = 16'h10a2; 14'h37ea: x = 16'h10a1; 14'h37eb: x = 16'h10a0; 14'h37ec: x = 16'h109f; 14'h37ed: x = 16'h109e; 14'h37ee: x = 16'h109d; 14'h37ef: x = 16'h109c; 14'h37f0: x = 16'h109b; 14'h37f1: x = 16'h109a; 14'h37f2: x = 16'h1098; 14'h37f3: x = 16'h1097; 14'h37f4: x = 16'h1096; 14'h37f5: x = 16'h1095; 14'h37f6: x = 16'h1094; 14'h37f7: x = 16'h1093; 14'h37f8: x = 16'h1092; 14'h37f9: x = 16'h1091; 14'h37fa: x = 16'h1090; 14'h37fb: x = 16'h108e; 14'h37fc: x = 16'h108d; 14'h37fd: x = 16'h108c; 14'h37fe: x = 16'h108b; 14'h37ff: x = 16'h108a; 14'h3800: x = 16'h1089; 14'h3801: x = 16'h1088; 14'h3802: x = 16'h1087; 14'h3803: x = 16'h1086; 14'h3804: x = 16'h1085; 14'h3805: x = 16'h1083; 14'h3806: x = 16'h1082; 14'h3807: x = 16'h1081; 14'h3808: x = 16'h1080; 14'h3809: x = 16'h107f; 14'h380a: x = 16'h107e; 14'h380b: x = 16'h107d; 14'h380c: x = 16'h107c; 14'h380d: x = 16'h107b; 14'h380e: x = 16'h1079; 14'h380f: x = 16'h1078; 14'h3810: x = 16'h1077; 14'h3811: x = 16'h1076; 14'h3812: x = 16'h1075; 14'h3813: x = 16'h1074; 14'h3814: x = 16'h1073; 14'h3815: x = 16'h1072; 14'h3816: x = 16'h1071; 14'h3817: x = 16'h106f; 14'h3818: x = 16'h106e; 14'h3819: x = 16'h106d; 14'h381a: x = 16'h106c; 14'h381b: x = 16'h106b; 14'h381c: x = 16'h106a; 14'h381d: x = 16'h1069; 14'h381e: x = 16'h1068; 14'h381f: x = 16'h1067; 14'h3820: x = 16'h1065; 14'h3821: x = 16'h1064; 14'h3822: x = 16'h1063; 14'h3823: x = 16'h1062; 14'h3824: x = 16'h1061; 14'h3825: x = 16'h1060; 14'h3826: x = 16'h105f; 14'h3827: x = 16'h105e; 14'h3828: x = 16'h105d; 14'h3829: x = 16'h105b; 14'h382a: x = 16'h105a; 14'h382b: x = 16'h1059; 14'h382c: x = 16'h1058; 14'h382d: x = 16'h1057; 14'h382e: x = 16'h1056; 14'h382f: x = 16'h1055; 14'h3830: x = 16'h1054; 14'h3831: x = 16'h1053; 14'h3832: x = 16'h1051; 14'h3833: x = 16'h1050; 14'h3834: x = 16'h104f; 14'h3835: x = 16'h104e; 14'h3836: x = 16'h104d; 14'h3837: x = 16'h104c; 14'h3838: x = 16'h104b; 14'h3839: x = 16'h104a; 14'h383a: x = 16'h1048; 14'h383b: x = 16'h1047; 14'h383c: x = 16'h1046; 14'h383d: x = 16'h1045; 14'h383e: x = 16'h1044; 14'h383f: x = 16'h1043; 14'h3840: x = 16'h1042; 14'h3841: x = 16'h1041; 14'h3842: x = 16'h1040; 14'h3843: x = 16'h103e; 14'h3844: x = 16'h103d; 14'h3845: x = 16'h103c; 14'h3846: x = 16'h103b; 14'h3847: x = 16'h103a; 14'h3848: x = 16'h1039; 14'h3849: x = 16'h1038; 14'h384a: x = 16'h1037; 14'h384b: x = 16'h1035; 14'h384c: x = 16'h1034; 14'h384d: x = 16'h1033; 14'h384e: x = 16'h1032; 14'h384f: x = 16'h1031; 14'h3850: x = 16'h1030; 14'h3851: x = 16'h102f; 14'h3852: x = 16'h102e; 14'h3853: x = 16'h102c; 14'h3854: x = 16'h102b; 14'h3855: x = 16'h102a; 14'h3856: x = 16'h1029; 14'h3857: x = 16'h1028; 14'h3858: x = 16'h1027; 14'h3859: x = 16'h1026; 14'h385a: x = 16'h1025; 14'h385b: x = 16'h1023; 14'h385c: x = 16'h1022; 14'h385d: x = 16'h1021; 14'h385e: x = 16'h1020; 14'h385f: x = 16'h101f; 14'h3860: x = 16'h101e; 14'h3861: x = 16'h101d; 14'h3862: x = 16'h101c; 14'h3863: x = 16'h101a; 14'h3864: x = 16'h1019; 14'h3865: x = 16'h1018; 14'h3866: x = 16'h1017; 14'h3867: x = 16'h1016; 14'h3868: x = 16'h1015; 14'h3869: x = 16'h1014; 14'h386a: x = 16'h1013; 14'h386b: x = 16'h1011; 14'h386c: x = 16'h1010; 14'h386d: x = 16'h100f; 14'h386e: x = 16'h100e; 14'h386f: x = 16'h100d; 14'h3870: x = 16'h100c; 14'h3871: x = 16'h100b; 14'h3872: x = 16'h1009; 14'h3873: x = 16'h1008; 14'h3874: x = 16'h1007; 14'h3875: x = 16'h1006; 14'h3876: x = 16'h1005; 14'h3877: x = 16'h1004; 14'h3878: x = 16'h1003; 14'h3879: x = 16'h1002; 14'h387a: x = 16'h1000; 14'h387b: x = 16'h fff; 14'h387c: x = 16'h ffe; 14'h387d: x = 16'h ffd; 14'h387e: x = 16'h ffc; 14'h387f: x = 16'h ffb; 14'h3880: x = 16'h ffa; 14'h3881: x = 16'h ff9; 14'h3882: x = 16'h ff7; 14'h3883: x = 16'h ff6; 14'h3884: x = 16'h ff5; 14'h3885: x = 16'h ff4; 14'h3886: x = 16'h ff3; 14'h3887: x = 16'h ff2; 14'h3888: x = 16'h ff1; 14'h3889: x = 16'h fef; 14'h388a: x = 16'h fee; 14'h388b: x = 16'h fed; 14'h388c: x = 16'h fec; 14'h388d: x = 16'h feb; 14'h388e: x = 16'h fea; 14'h388f: x = 16'h fe9; 14'h3890: x = 16'h fe7; 14'h3891: x = 16'h fe6; 14'h3892: x = 16'h fe5; 14'h3893: x = 16'h fe4; 14'h3894: x = 16'h fe3; 14'h3895: x = 16'h fe2; 14'h3896: x = 16'h fe1; 14'h3897: x = 16'h fdf; 14'h3898: x = 16'h fde; 14'h3899: x = 16'h fdd; 14'h389a: x = 16'h fdc; 14'h389b: x = 16'h fdb; 14'h389c: x = 16'h fda; 14'h389d: x = 16'h fd9; 14'h389e: x = 16'h fd7; 14'h389f: x = 16'h fd6; 14'h38a0: x = 16'h fd5; 14'h38a1: x = 16'h fd4; 14'h38a2: x = 16'h fd3; 14'h38a3: x = 16'h fd2; 14'h38a4: x = 16'h fd1; 14'h38a5: x = 16'h fd0; 14'h38a6: x = 16'h fce; 14'h38a7: x = 16'h fcd; 14'h38a8: x = 16'h fcc; 14'h38a9: x = 16'h fcb; 14'h38aa: x = 16'h fca; 14'h38ab: x = 16'h fc9; 14'h38ac: x = 16'h fc7; 14'h38ad: x = 16'h fc6; 14'h38ae: x = 16'h fc5; 14'h38af: x = 16'h fc4; 14'h38b0: x = 16'h fc3; 14'h38b1: x = 16'h fc2; 14'h38b2: x = 16'h fc1; 14'h38b3: x = 16'h fbf; 14'h38b4: x = 16'h fbe; 14'h38b5: x = 16'h fbd; 14'h38b6: x = 16'h fbc; 14'h38b7: x = 16'h fbb; 14'h38b8: x = 16'h fba; 14'h38b9: x = 16'h fb9; 14'h38ba: x = 16'h fb7; 14'h38bb: x = 16'h fb6; 14'h38bc: x = 16'h fb5; 14'h38bd: x = 16'h fb4; 14'h38be: x = 16'h fb3; 14'h38bf: x = 16'h fb2; 14'h38c0: x = 16'h fb1; 14'h38c1: x = 16'h faf; 14'h38c2: x = 16'h fae; 14'h38c3: x = 16'h fad; 14'h38c4: x = 16'h fac; 14'h38c5: x = 16'h fab; 14'h38c6: x = 16'h faa; 14'h38c7: x = 16'h fa8; 14'h38c8: x = 16'h fa7; 14'h38c9: x = 16'h fa6; 14'h38ca: x = 16'h fa5; 14'h38cb: x = 16'h fa4; 14'h38cc: x = 16'h fa3; 14'h38cd: x = 16'h fa2; 14'h38ce: x = 16'h fa0; 14'h38cf: x = 16'h f9f; 14'h38d0: x = 16'h f9e; 14'h38d1: x = 16'h f9d; 14'h38d2: x = 16'h f9c; 14'h38d3: x = 16'h f9b; 14'h38d4: x = 16'h f99; 14'h38d5: x = 16'h f98; 14'h38d6: x = 16'h f97; 14'h38d7: x = 16'h f96; 14'h38d8: x = 16'h f95; 14'h38d9: x = 16'h f94; 14'h38da: x = 16'h f93; 14'h38db: x = 16'h f91; 14'h38dc: x = 16'h f90; 14'h38dd: x = 16'h f8f; 14'h38de: x = 16'h f8e; 14'h38df: x = 16'h f8d; 14'h38e0: x = 16'h f8c; 14'h38e1: x = 16'h f8a; 14'h38e2: x = 16'h f89; 14'h38e3: x = 16'h f88; 14'h38e4: x = 16'h f87; 14'h38e5: x = 16'h f86; 14'h38e6: x = 16'h f85; 14'h38e7: x = 16'h f84; 14'h38e8: x = 16'h f82; 14'h38e9: x = 16'h f81; 14'h38ea: x = 16'h f80; 14'h38eb: x = 16'h f7f; 14'h38ec: x = 16'h f7e; 14'h38ed: x = 16'h f7d; 14'h38ee: x = 16'h f7b; 14'h38ef: x = 16'h f7a; 14'h38f0: x = 16'h f79; 14'h38f1: x = 16'h f78; 14'h38f2: x = 16'h f77; 14'h38f3: x = 16'h f76; 14'h38f4: x = 16'h f74; 14'h38f5: x = 16'h f73; 14'h38f6: x = 16'h f72; 14'h38f7: x = 16'h f71; 14'h38f8: x = 16'h f70; 14'h38f9: x = 16'h f6f; 14'h38fa: x = 16'h f6d; 14'h38fb: x = 16'h f6c; 14'h38fc: x = 16'h f6b; 14'h38fd: x = 16'h f6a; 14'h38fe: x = 16'h f69; 14'h38ff: x = 16'h f68; 14'h3900: x = 16'h f66; 14'h3901: x = 16'h f65; 14'h3902: x = 16'h f64; 14'h3903: x = 16'h f63; 14'h3904: x = 16'h f62; 14'h3905: x = 16'h f61; 14'h3906: x = 16'h f5f; 14'h3907: x = 16'h f5e; 14'h3908: x = 16'h f5d; 14'h3909: x = 16'h f5c; 14'h390a: x = 16'h f5b; 14'h390b: x = 16'h f5a; 14'h390c: x = 16'h f58; 14'h390d: x = 16'h f57; 14'h390e: x = 16'h f56; 14'h390f: x = 16'h f55; 14'h3910: x = 16'h f54; 14'h3911: x = 16'h f53; 14'h3912: x = 16'h f51; 14'h3913: x = 16'h f50; 14'h3914: x = 16'h f4f; 14'h3915: x = 16'h f4e; 14'h3916: x = 16'h f4d; 14'h3917: x = 16'h f4c; 14'h3918: x = 16'h f4a; 14'h3919: x = 16'h f49; 14'h391a: x = 16'h f48; 14'h391b: x = 16'h f47; 14'h391c: x = 16'h f46; 14'h391d: x = 16'h f44; 14'h391e: x = 16'h f43; 14'h391f: x = 16'h f42; 14'h3920: x = 16'h f41; 14'h3921: x = 16'h f40; 14'h3922: x = 16'h f3f; 14'h3923: x = 16'h f3d; 14'h3924: x = 16'h f3c; 14'h3925: x = 16'h f3b; 14'h3926: x = 16'h f3a; 14'h3927: x = 16'h f39; 14'h3928: x = 16'h f38; 14'h3929: x = 16'h f36; 14'h392a: x = 16'h f35; 14'h392b: x = 16'h f34; 14'h392c: x = 16'h f33; 14'h392d: x = 16'h f32; 14'h392e: x = 16'h f30; 14'h392f: x = 16'h f2f; 14'h3930: x = 16'h f2e; 14'h3931: x = 16'h f2d; 14'h3932: x = 16'h f2c; 14'h3933: x = 16'h f2b; 14'h3934: x = 16'h f29; 14'h3935: x = 16'h f28; 14'h3936: x = 16'h f27; 14'h3937: x = 16'h f26; 14'h3938: x = 16'h f25; 14'h3939: x = 16'h f24; 14'h393a: x = 16'h f22; 14'h393b: x = 16'h f21; 14'h393c: x = 16'h f20; 14'h393d: x = 16'h f1f; 14'h393e: x = 16'h f1e; 14'h393f: x = 16'h f1c; 14'h3940: x = 16'h f1b; 14'h3941: x = 16'h f1a; 14'h3942: x = 16'h f19; 14'h3943: x = 16'h f18; 14'h3944: x = 16'h f16; 14'h3945: x = 16'h f15; 14'h3946: x = 16'h f14; 14'h3947: x = 16'h f13; 14'h3948: x = 16'h f12; 14'h3949: x = 16'h f11; 14'h394a: x = 16'h f0f; 14'h394b: x = 16'h f0e; 14'h394c: x = 16'h f0d; 14'h394d: x = 16'h f0c; 14'h394e: x = 16'h f0b; 14'h394f: x = 16'h f09; 14'h3950: x = 16'h f08; 14'h3951: x = 16'h f07; 14'h3952: x = 16'h f06; 14'h3953: x = 16'h f05; 14'h3954: x = 16'h f03; 14'h3955: x = 16'h f02; 14'h3956: x = 16'h f01; 14'h3957: x = 16'h f00; 14'h3958: x = 16'h eff; 14'h3959: x = 16'h efe; 14'h395a: x = 16'h efc; 14'h395b: x = 16'h efb; 14'h395c: x = 16'h efa; 14'h395d: x = 16'h ef9; 14'h395e: x = 16'h ef8; 14'h395f: x = 16'h ef6; 14'h3960: x = 16'h ef5; 14'h3961: x = 16'h ef4; 14'h3962: x = 16'h ef3; 14'h3963: x = 16'h ef2; 14'h3964: x = 16'h ef0; 14'h3965: x = 16'h eef; 14'h3966: x = 16'h eee; 14'h3967: x = 16'h eed; 14'h3968: x = 16'h eec; 14'h3969: x = 16'h eea; 14'h396a: x = 16'h ee9; 14'h396b: x = 16'h ee8; 14'h396c: x = 16'h ee7; 14'h396d: x = 16'h ee6; 14'h396e: x = 16'h ee4; 14'h396f: x = 16'h ee3; 14'h3970: x = 16'h ee2; 14'h3971: x = 16'h ee1; 14'h3972: x = 16'h ee0; 14'h3973: x = 16'h ede; 14'h3974: x = 16'h edd; 14'h3975: x = 16'h edc; 14'h3976: x = 16'h edb; 14'h3977: x = 16'h eda; 14'h3978: x = 16'h ed8; 14'h3979: x = 16'h ed7; 14'h397a: x = 16'h ed6; 14'h397b: x = 16'h ed5; 14'h397c: x = 16'h ed4; 14'h397d: x = 16'h ed2; 14'h397e: x = 16'h ed1; 14'h397f: x = 16'h ed0; 14'h3980: x = 16'h ecf; 14'h3981: x = 16'h ece; 14'h3982: x = 16'h ecc; 14'h3983: x = 16'h ecb; 14'h3984: x = 16'h eca; 14'h3985: x = 16'h ec9; 14'h3986: x = 16'h ec8; 14'h3987: x = 16'h ec6; 14'h3988: x = 16'h ec5; 14'h3989: x = 16'h ec4; 14'h398a: x = 16'h ec3; 14'h398b: x = 16'h ec2; 14'h398c: x = 16'h ec0; 14'h398d: x = 16'h ebf; 14'h398e: x = 16'h ebe; 14'h398f: x = 16'h ebd; 14'h3990: x = 16'h ebc; 14'h3991: x = 16'h eba; 14'h3992: x = 16'h eb9; 14'h3993: x = 16'h eb8; 14'h3994: x = 16'h eb7; 14'h3995: x = 16'h eb6; 14'h3996: x = 16'h eb4; 14'h3997: x = 16'h eb3; 14'h3998: x = 16'h eb2; 14'h3999: x = 16'h eb1; 14'h399a: x = 16'h eb0; 14'h399b: x = 16'h eae; 14'h399c: x = 16'h ead; 14'h399d: x = 16'h eac; 14'h399e: x = 16'h eab; 14'h399f: x = 16'h ea9; 14'h39a0: x = 16'h ea8; 14'h39a1: x = 16'h ea7; 14'h39a2: x = 16'h ea6; 14'h39a3: x = 16'h ea5; 14'h39a4: x = 16'h ea3; 14'h39a5: x = 16'h ea2; 14'h39a6: x = 16'h ea1; 14'h39a7: x = 16'h ea0; 14'h39a8: x = 16'h e9f; 14'h39a9: x = 16'h e9d; 14'h39aa: x = 16'h e9c; 14'h39ab: x = 16'h e9b; 14'h39ac: x = 16'h e9a; 14'h39ad: x = 16'h e98; 14'h39ae: x = 16'h e97; 14'h39af: x = 16'h e96; 14'h39b0: x = 16'h e95; 14'h39b1: x = 16'h e94; 14'h39b2: x = 16'h e92; 14'h39b3: x = 16'h e91; 14'h39b4: x = 16'h e90; 14'h39b5: x = 16'h e8f; 14'h39b6: x = 16'h e8d; 14'h39b7: x = 16'h e8c; 14'h39b8: x = 16'h e8b; 14'h39b9: x = 16'h e8a; 14'h39ba: x = 16'h e89; 14'h39bb: x = 16'h e87; 14'h39bc: x = 16'h e86; 14'h39bd: x = 16'h e85; 14'h39be: x = 16'h e84; 14'h39bf: x = 16'h e83; 14'h39c0: x = 16'h e81; 14'h39c1: x = 16'h e80; 14'h39c2: x = 16'h e7f; 14'h39c3: x = 16'h e7e; 14'h39c4: x = 16'h e7c; 14'h39c5: x = 16'h e7b; 14'h39c6: x = 16'h e7a; 14'h39c7: x = 16'h e79; 14'h39c8: x = 16'h e77; 14'h39c9: x = 16'h e76; 14'h39ca: x = 16'h e75; 14'h39cb: x = 16'h e74; 14'h39cc: x = 16'h e73; 14'h39cd: x = 16'h e71; 14'h39ce: x = 16'h e70; 14'h39cf: x = 16'h e6f; 14'h39d0: x = 16'h e6e; 14'h39d1: x = 16'h e6c; 14'h39d2: x = 16'h e6b; 14'h39d3: x = 16'h e6a; 14'h39d4: x = 16'h e69; 14'h39d5: x = 16'h e68; 14'h39d6: x = 16'h e66; 14'h39d7: x = 16'h e65; 14'h39d8: x = 16'h e64; 14'h39d9: x = 16'h e63; 14'h39da: x = 16'h e61; 14'h39db: x = 16'h e60; 14'h39dc: x = 16'h e5f; 14'h39dd: x = 16'h e5e; 14'h39de: x = 16'h e5c; 14'h39df: x = 16'h e5b; 14'h39e0: x = 16'h e5a; 14'h39e1: x = 16'h e59; 14'h39e2: x = 16'h e58; 14'h39e3: x = 16'h e56; 14'h39e4: x = 16'h e55; 14'h39e5: x = 16'h e54; 14'h39e6: x = 16'h e53; 14'h39e7: x = 16'h e51; 14'h39e8: x = 16'h e50; 14'h39e9: x = 16'h e4f; 14'h39ea: x = 16'h e4e; 14'h39eb: x = 16'h e4c; 14'h39ec: x = 16'h e4b; 14'h39ed: x = 16'h e4a; 14'h39ee: x = 16'h e49; 14'h39ef: x = 16'h e47; 14'h39f0: x = 16'h e46; 14'h39f1: x = 16'h e45; 14'h39f2: x = 16'h e44; 14'h39f3: x = 16'h e43; 14'h39f4: x = 16'h e41; 14'h39f5: x = 16'h e40; 14'h39f6: x = 16'h e3f; 14'h39f7: x = 16'h e3e; 14'h39f8: x = 16'h e3c; 14'h39f9: x = 16'h e3b; 14'h39fa: x = 16'h e3a; 14'h39fb: x = 16'h e39; 14'h39fc: x = 16'h e37; 14'h39fd: x = 16'h e36; 14'h39fe: x = 16'h e35; 14'h39ff: x = 16'h e34; 14'h3a00: x = 16'h e32; 14'h3a01: x = 16'h e31; 14'h3a02: x = 16'h e30; 14'h3a03: x = 16'h e2f; 14'h3a04: x = 16'h e2d; 14'h3a05: x = 16'h e2c; 14'h3a06: x = 16'h e2b; 14'h3a07: x = 16'h e2a; 14'h3a08: x = 16'h e28; 14'h3a09: x = 16'h e27; 14'h3a0a: x = 16'h e26; 14'h3a0b: x = 16'h e25; 14'h3a0c: x = 16'h e23; 14'h3a0d: x = 16'h e22; 14'h3a0e: x = 16'h e21; 14'h3a0f: x = 16'h e20; 14'h3a10: x = 16'h e1e; 14'h3a11: x = 16'h e1d; 14'h3a12: x = 16'h e1c; 14'h3a13: x = 16'h e1b; 14'h3a14: x = 16'h e19; 14'h3a15: x = 16'h e18; 14'h3a16: x = 16'h e17; 14'h3a17: x = 16'h e16; 14'h3a18: x = 16'h e14; 14'h3a19: x = 16'h e13; 14'h3a1a: x = 16'h e12; 14'h3a1b: x = 16'h e11; 14'h3a1c: x = 16'h e0f; 14'h3a1d: x = 16'h e0e; 14'h3a1e: x = 16'h e0d; 14'h3a1f: x = 16'h e0c; 14'h3a20: x = 16'h e0a; 14'h3a21: x = 16'h e09; 14'h3a22: x = 16'h e08; 14'h3a23: x = 16'h e07; 14'h3a24: x = 16'h e05; 14'h3a25: x = 16'h e04; 14'h3a26: x = 16'h e03; 14'h3a27: x = 16'h e02; 14'h3a28: x = 16'h e00; 14'h3a29: x = 16'h dff; 14'h3a2a: x = 16'h dfe; 14'h3a2b: x = 16'h dfd; 14'h3a2c: x = 16'h dfb; 14'h3a2d: x = 16'h dfa; 14'h3a2e: x = 16'h df9; 14'h3a2f: x = 16'h df8; 14'h3a30: x = 16'h df6; 14'h3a31: x = 16'h df5; 14'h3a32: x = 16'h df4; 14'h3a33: x = 16'h df3; 14'h3a34: x = 16'h df1; 14'h3a35: x = 16'h df0; 14'h3a36: x = 16'h def; 14'h3a37: x = 16'h ded; 14'h3a38: x = 16'h dec; 14'h3a39: x = 16'h deb; 14'h3a3a: x = 16'h dea; 14'h3a3b: x = 16'h de8; 14'h3a3c: x = 16'h de7; 14'h3a3d: x = 16'h de6; 14'h3a3e: x = 16'h de5; 14'h3a3f: x = 16'h de3; 14'h3a40: x = 16'h de2; 14'h3a41: x = 16'h de1; 14'h3a42: x = 16'h de0; 14'h3a43: x = 16'h dde; 14'h3a44: x = 16'h ddd; 14'h3a45: x = 16'h ddc; 14'h3a46: x = 16'h dda; 14'h3a47: x = 16'h dd9; 14'h3a48: x = 16'h dd8; 14'h3a49: x = 16'h dd7; 14'h3a4a: x = 16'h dd5; 14'h3a4b: x = 16'h dd4; 14'h3a4c: x = 16'h dd3; 14'h3a4d: x = 16'h dd2; 14'h3a4e: x = 16'h dd0; 14'h3a4f: x = 16'h dcf; 14'h3a50: x = 16'h dce; 14'h3a51: x = 16'h dcd; 14'h3a52: x = 16'h dcb; 14'h3a53: x = 16'h dca; 14'h3a54: x = 16'h dc9; 14'h3a55: x = 16'h dc7; 14'h3a56: x = 16'h dc6; 14'h3a57: x = 16'h dc5; 14'h3a58: x = 16'h dc4; 14'h3a59: x = 16'h dc2; 14'h3a5a: x = 16'h dc1; 14'h3a5b: x = 16'h dc0; 14'h3a5c: x = 16'h dbe; 14'h3a5d: x = 16'h dbd; 14'h3a5e: x = 16'h dbc; 14'h3a5f: x = 16'h dbb; 14'h3a60: x = 16'h db9; 14'h3a61: x = 16'h db8; 14'h3a62: x = 16'h db7; 14'h3a63: x = 16'h db6; 14'h3a64: x = 16'h db4; 14'h3a65: x = 16'h db3; 14'h3a66: x = 16'h db2; 14'h3a67: x = 16'h db0; 14'h3a68: x = 16'h daf; 14'h3a69: x = 16'h dae; 14'h3a6a: x = 16'h dad; 14'h3a6b: x = 16'h dab; 14'h3a6c: x = 16'h daa; 14'h3a6d: x = 16'h da9; 14'h3a6e: x = 16'h da7; 14'h3a6f: x = 16'h da6; 14'h3a70: x = 16'h da5; 14'h3a71: x = 16'h da4; 14'h3a72: x = 16'h da2; 14'h3a73: x = 16'h da1; 14'h3a74: x = 16'h da0; 14'h3a75: x = 16'h d9e; 14'h3a76: x = 16'h d9d; 14'h3a77: x = 16'h d9c; 14'h3a78: x = 16'h d9b; 14'h3a79: x = 16'h d99; 14'h3a7a: x = 16'h d98; 14'h3a7b: x = 16'h d97; 14'h3a7c: x = 16'h d95; 14'h3a7d: x = 16'h d94; 14'h3a7e: x = 16'h d93; 14'h3a7f: x = 16'h d92; 14'h3a80: x = 16'h d90; 14'h3a81: x = 16'h d8f; 14'h3a82: x = 16'h d8e; 14'h3a83: x = 16'h d8c; 14'h3a84: x = 16'h d8b; 14'h3a85: x = 16'h d8a; 14'h3a86: x = 16'h d89; 14'h3a87: x = 16'h d87; 14'h3a88: x = 16'h d86; 14'h3a89: x = 16'h d85; 14'h3a8a: x = 16'h d83; 14'h3a8b: x = 16'h d82; 14'h3a8c: x = 16'h d81; 14'h3a8d: x = 16'h d7f; 14'h3a8e: x = 16'h d7e; 14'h3a8f: x = 16'h d7d; 14'h3a90: x = 16'h d7c; 14'h3a91: x = 16'h d7a; 14'h3a92: x = 16'h d79; 14'h3a93: x = 16'h d78; 14'h3a94: x = 16'h d76; 14'h3a95: x = 16'h d75; 14'h3a96: x = 16'h d74; 14'h3a97: x = 16'h d73; 14'h3a98: x = 16'h d71; 14'h3a99: x = 16'h d70; 14'h3a9a: x = 16'h d6f; 14'h3a9b: x = 16'h d6d; 14'h3a9c: x = 16'h d6c; 14'h3a9d: x = 16'h d6b; 14'h3a9e: x = 16'h d69; 14'h3a9f: x = 16'h d68; 14'h3aa0: x = 16'h d67; 14'h3aa1: x = 16'h d65; 14'h3aa2: x = 16'h d64; 14'h3aa3: x = 16'h d63; 14'h3aa4: x = 16'h d62; 14'h3aa5: x = 16'h d60; 14'h3aa6: x = 16'h d5f; 14'h3aa7: x = 16'h d5e; 14'h3aa8: x = 16'h d5c; 14'h3aa9: x = 16'h d5b; 14'h3aaa: x = 16'h d5a; 14'h3aab: x = 16'h d58; 14'h3aac: x = 16'h d57; 14'h3aad: x = 16'h d56; 14'h3aae: x = 16'h d55; 14'h3aaf: x = 16'h d53; 14'h3ab0: x = 16'h d52; 14'h3ab1: x = 16'h d51; 14'h3ab2: x = 16'h d4f; 14'h3ab3: x = 16'h d4e; 14'h3ab4: x = 16'h d4d; 14'h3ab5: x = 16'h d4b; 14'h3ab6: x = 16'h d4a; 14'h3ab7: x = 16'h d49; 14'h3ab8: x = 16'h d47; 14'h3ab9: x = 16'h d46; 14'h3aba: x = 16'h d45; 14'h3abb: x = 16'h d43; 14'h3abc: x = 16'h d42; 14'h3abd: x = 16'h d41; 14'h3abe: x = 16'h d40; 14'h3abf: x = 16'h d3e; 14'h3ac0: x = 16'h d3d; 14'h3ac1: x = 16'h d3c; 14'h3ac2: x = 16'h d3a; 14'h3ac3: x = 16'h d39; 14'h3ac4: x = 16'h d38; 14'h3ac5: x = 16'h d36; 14'h3ac6: x = 16'h d35; 14'h3ac7: x = 16'h d34; 14'h3ac8: x = 16'h d32; 14'h3ac9: x = 16'h d31; 14'h3aca: x = 16'h d30; 14'h3acb: x = 16'h d2e; 14'h3acc: x = 16'h d2d; 14'h3acd: x = 16'h d2c; 14'h3ace: x = 16'h d2a; 14'h3acf: x = 16'h d29; 14'h3ad0: x = 16'h d28; 14'h3ad1: x = 16'h d26; 14'h3ad2: x = 16'h d25; 14'h3ad3: x = 16'h d24; 14'h3ad4: x = 16'h d22; 14'h3ad5: x = 16'h d21; 14'h3ad6: x = 16'h d20; 14'h3ad7: x = 16'h d1e; 14'h3ad8: x = 16'h d1d; 14'h3ad9: x = 16'h d1c; 14'h3ada: x = 16'h d1b; 14'h3adb: x = 16'h d19; 14'h3adc: x = 16'h d18; 14'h3add: x = 16'h d17; 14'h3ade: x = 16'h d15; 14'h3adf: x = 16'h d14; 14'h3ae0: x = 16'h d13; 14'h3ae1: x = 16'h d11; 14'h3ae2: x = 16'h d10; 14'h3ae3: x = 16'h d0f; 14'h3ae4: x = 16'h d0d; 14'h3ae5: x = 16'h d0c; 14'h3ae6: x = 16'h d0b; 14'h3ae7: x = 16'h d09; 14'h3ae8: x = 16'h d08; 14'h3ae9: x = 16'h d07; 14'h3aea: x = 16'h d05; 14'h3aeb: x = 16'h d04; 14'h3aec: x = 16'h d03; 14'h3aed: x = 16'h d01; 14'h3aee: x = 16'h d00; 14'h3aef: x = 16'h cff; 14'h3af0: x = 16'h cfd; 14'h3af1: x = 16'h cfc; 14'h3af2: x = 16'h cfb; 14'h3af3: x = 16'h cf9; 14'h3af4: x = 16'h cf8; 14'h3af5: x = 16'h cf7; 14'h3af6: x = 16'h cf5; 14'h3af7: x = 16'h cf4; 14'h3af8: x = 16'h cf2; 14'h3af9: x = 16'h cf1; 14'h3afa: x = 16'h cf0; 14'h3afb: x = 16'h cee; 14'h3afc: x = 16'h ced; 14'h3afd: x = 16'h cec; 14'h3afe: x = 16'h cea; 14'h3aff: x = 16'h ce9; 14'h3b00: x = 16'h ce8; 14'h3b01: x = 16'h ce6; 14'h3b02: x = 16'h ce5; 14'h3b03: x = 16'h ce4; 14'h3b04: x = 16'h ce2; 14'h3b05: x = 16'h ce1; 14'h3b06: x = 16'h ce0; 14'h3b07: x = 16'h cde; 14'h3b08: x = 16'h cdd; 14'h3b09: x = 16'h cdc; 14'h3b0a: x = 16'h cda; 14'h3b0b: x = 16'h cd9; 14'h3b0c: x = 16'h cd8; 14'h3b0d: x = 16'h cd6; 14'h3b0e: x = 16'h cd5; 14'h3b0f: x = 16'h cd4; 14'h3b10: x = 16'h cd2; 14'h3b11: x = 16'h cd1; 14'h3b12: x = 16'h ccf; 14'h3b13: x = 16'h cce; 14'h3b14: x = 16'h ccd; 14'h3b15: x = 16'h ccb; 14'h3b16: x = 16'h cca; 14'h3b17: x = 16'h cc9; 14'h3b18: x = 16'h cc7; 14'h3b19: x = 16'h cc6; 14'h3b1a: x = 16'h cc5; 14'h3b1b: x = 16'h cc3; 14'h3b1c: x = 16'h cc2; 14'h3b1d: x = 16'h cc1; 14'h3b1e: x = 16'h cbf; 14'h3b1f: x = 16'h cbe; 14'h3b20: x = 16'h cbc; 14'h3b21: x = 16'h cbb; 14'h3b22: x = 16'h cba; 14'h3b23: x = 16'h cb8; 14'h3b24: x = 16'h cb7; 14'h3b25: x = 16'h cb6; 14'h3b26: x = 16'h cb4; 14'h3b27: x = 16'h cb3; 14'h3b28: x = 16'h cb2; 14'h3b29: x = 16'h cb0; 14'h3b2a: x = 16'h caf; 14'h3b2b: x = 16'h cad; 14'h3b2c: x = 16'h cac; 14'h3b2d: x = 16'h cab; 14'h3b2e: x = 16'h ca9; 14'h3b2f: x = 16'h ca8; 14'h3b30: x = 16'h ca7; 14'h3b31: x = 16'h ca5; 14'h3b32: x = 16'h ca4; 14'h3b33: x = 16'h ca3; 14'h3b34: x = 16'h ca1; 14'h3b35: x = 16'h ca0; 14'h3b36: x = 16'h c9e; 14'h3b37: x = 16'h c9d; 14'h3b38: x = 16'h c9c; 14'h3b39: x = 16'h c9a; 14'h3b3a: x = 16'h c99; 14'h3b3b: x = 16'h c98; 14'h3b3c: x = 16'h c96; 14'h3b3d: x = 16'h c95; 14'h3b3e: x = 16'h c93; 14'h3b3f: x = 16'h c92; 14'h3b40: x = 16'h c91; 14'h3b41: x = 16'h c8f; 14'h3b42: x = 16'h c8e; 14'h3b43: x = 16'h c8d; 14'h3b44: x = 16'h c8b; 14'h3b45: x = 16'h c8a; 14'h3b46: x = 16'h c88; 14'h3b47: x = 16'h c87; 14'h3b48: x = 16'h c86; 14'h3b49: x = 16'h c84; 14'h3b4a: x = 16'h c83; 14'h3b4b: x = 16'h c82; 14'h3b4c: x = 16'h c80; 14'h3b4d: x = 16'h c7f; 14'h3b4e: x = 16'h c7d; 14'h3b4f: x = 16'h c7c; 14'h3b50: x = 16'h c7b; 14'h3b51: x = 16'h c79; 14'h3b52: x = 16'h c78; 14'h3b53: x = 16'h c77; 14'h3b54: x = 16'h c75; 14'h3b55: x = 16'h c74; 14'h3b56: x = 16'h c72; 14'h3b57: x = 16'h c71; 14'h3b58: x = 16'h c70; 14'h3b59: x = 16'h c6e; 14'h3b5a: x = 16'h c6d; 14'h3b5b: x = 16'h c6b; 14'h3b5c: x = 16'h c6a; 14'h3b5d: x = 16'h c69; 14'h3b5e: x = 16'h c67; 14'h3b5f: x = 16'h c66; 14'h3b60: x = 16'h c64; 14'h3b61: x = 16'h c63; 14'h3b62: x = 16'h c62; 14'h3b63: x = 16'h c60; 14'h3b64: x = 16'h c5f; 14'h3b65: x = 16'h c5d; 14'h3b66: x = 16'h c5c; 14'h3b67: x = 16'h c5b; 14'h3b68: x = 16'h c59; 14'h3b69: x = 16'h c58; 14'h3b6a: x = 16'h c57; 14'h3b6b: x = 16'h c55; 14'h3b6c: x = 16'h c54; 14'h3b6d: x = 16'h c52; 14'h3b6e: x = 16'h c51; 14'h3b6f: x = 16'h c50; 14'h3b70: x = 16'h c4e; 14'h3b71: x = 16'h c4d; 14'h3b72: x = 16'h c4b; 14'h3b73: x = 16'h c4a; 14'h3b74: x = 16'h c49; 14'h3b75: x = 16'h c47; 14'h3b76: x = 16'h c46; 14'h3b77: x = 16'h c44; 14'h3b78: x = 16'h c43; 14'h3b79: x = 16'h c42; 14'h3b7a: x = 16'h c40; 14'h3b7b: x = 16'h c3f; 14'h3b7c: x = 16'h c3d; 14'h3b7d: x = 16'h c3c; 14'h3b7e: x = 16'h c3a; 14'h3b7f: x = 16'h c39; 14'h3b80: x = 16'h c38; 14'h3b81: x = 16'h c36; 14'h3b82: x = 16'h c35; 14'h3b83: x = 16'h c33; 14'h3b84: x = 16'h c32; 14'h3b85: x = 16'h c31; 14'h3b86: x = 16'h c2f; 14'h3b87: x = 16'h c2e; 14'h3b88: x = 16'h c2c; 14'h3b89: x = 16'h c2b; 14'h3b8a: x = 16'h c2a; 14'h3b8b: x = 16'h c28; 14'h3b8c: x = 16'h c27; 14'h3b8d: x = 16'h c25; 14'h3b8e: x = 16'h c24; 14'h3b8f: x = 16'h c22; 14'h3b90: x = 16'h c21; 14'h3b91: x = 16'h c20; 14'h3b92: x = 16'h c1e; 14'h3b93: x = 16'h c1d; 14'h3b94: x = 16'h c1b; 14'h3b95: x = 16'h c1a; 14'h3b96: x = 16'h c19; 14'h3b97: x = 16'h c17; 14'h3b98: x = 16'h c16; 14'h3b99: x = 16'h c14; 14'h3b9a: x = 16'h c13; 14'h3b9b: x = 16'h c11; 14'h3b9c: x = 16'h c10; 14'h3b9d: x = 16'h c0f; 14'h3b9e: x = 16'h c0d; 14'h3b9f: x = 16'h c0c; 14'h3ba0: x = 16'h c0a; 14'h3ba1: x = 16'h c09; 14'h3ba2: x = 16'h c07; 14'h3ba3: x = 16'h c06; 14'h3ba4: x = 16'h c05; 14'h3ba5: x = 16'h c03; 14'h3ba6: x = 16'h c02; 14'h3ba7: x = 16'h c00; 14'h3ba8: x = 16'h bff; 14'h3ba9: x = 16'h bfd; 14'h3baa: x = 16'h bfc; 14'h3bab: x = 16'h bfb; 14'h3bac: x = 16'h bf9; 14'h3bad: x = 16'h bf8; 14'h3bae: x = 16'h bf6; 14'h3baf: x = 16'h bf5; 14'h3bb0: x = 16'h bf3; 14'h3bb1: x = 16'h bf2; 14'h3bb2: x = 16'h bf1; 14'h3bb3: x = 16'h bef; 14'h3bb4: x = 16'h bee; 14'h3bb5: x = 16'h bec; 14'h3bb6: x = 16'h beb; 14'h3bb7: x = 16'h be9; 14'h3bb8: x = 16'h be8; 14'h3bb9: x = 16'h be6; 14'h3bba: x = 16'h be5; 14'h3bbb: x = 16'h be4; 14'h3bbc: x = 16'h be2; 14'h3bbd: x = 16'h be1; 14'h3bbe: x = 16'h bdf; 14'h3bbf: x = 16'h bde; 14'h3bc0: x = 16'h bdc; 14'h3bc1: x = 16'h bdb; 14'h3bc2: x = 16'h bd9; 14'h3bc3: x = 16'h bd8; 14'h3bc4: x = 16'h bd7; 14'h3bc5: x = 16'h bd5; 14'h3bc6: x = 16'h bd4; 14'h3bc7: x = 16'h bd2; 14'h3bc8: x = 16'h bd1; 14'h3bc9: x = 16'h bcf; 14'h3bca: x = 16'h bce; 14'h3bcb: x = 16'h bcc; 14'h3bcc: x = 16'h bcb; 14'h3bcd: x = 16'h bca; 14'h3bce: x = 16'h bc8; 14'h3bcf: x = 16'h bc7; 14'h3bd0: x = 16'h bc5; 14'h3bd1: x = 16'h bc4; 14'h3bd2: x = 16'h bc2; 14'h3bd3: x = 16'h bc1; 14'h3bd4: x = 16'h bbf; 14'h3bd5: x = 16'h bbe; 14'h3bd6: x = 16'h bbc; 14'h3bd7: x = 16'h bbb; 14'h3bd8: x = 16'h bba; 14'h3bd9: x = 16'h bb8; 14'h3bda: x = 16'h bb7; 14'h3bdb: x = 16'h bb5; 14'h3bdc: x = 16'h bb4; 14'h3bdd: x = 16'h bb2; 14'h3bde: x = 16'h bb1; 14'h3bdf: x = 16'h baf; 14'h3be0: x = 16'h bae; 14'h3be1: x = 16'h bac; 14'h3be2: x = 16'h bab; 14'h3be3: x = 16'h ba9; 14'h3be4: x = 16'h ba8; 14'h3be5: x = 16'h ba7; 14'h3be6: x = 16'h ba5; 14'h3be7: x = 16'h ba4; 14'h3be8: x = 16'h ba2; 14'h3be9: x = 16'h ba1; 14'h3bea: x = 16'h b9f; 14'h3beb: x = 16'h b9e; 14'h3bec: x = 16'h b9c; 14'h3bed: x = 16'h b9b; 14'h3bee: x = 16'h b99; 14'h3bef: x = 16'h b98; 14'h3bf0: x = 16'h b96; 14'h3bf1: x = 16'h b95; 14'h3bf2: x = 16'h b93; 14'h3bf3: x = 16'h b92; 14'h3bf4: x = 16'h b90; 14'h3bf5: x = 16'h b8f; 14'h3bf6: x = 16'h b8d; 14'h3bf7: x = 16'h b8c; 14'h3bf8: x = 16'h b8b; 14'h3bf9: x = 16'h b89; 14'h3bfa: x = 16'h b88; 14'h3bfb: x = 16'h b86; 14'h3bfc: x = 16'h b85; 14'h3bfd: x = 16'h b83; 14'h3bfe: x = 16'h b82; 14'h3bff: x = 16'h b80; 14'h3c00: x = 16'h b7f; 14'h3c01: x = 16'h b7d; 14'h3c02: x = 16'h b7c; 14'h3c03: x = 16'h b7a; 14'h3c04: x = 16'h b79; 14'h3c05: x = 16'h b77; 14'h3c06: x = 16'h b76; 14'h3c07: x = 16'h b74; 14'h3c08: x = 16'h b73; 14'h3c09: x = 16'h b71; 14'h3c0a: x = 16'h b70; 14'h3c0b: x = 16'h b6e; 14'h3c0c: x = 16'h b6d; 14'h3c0d: x = 16'h b6b; 14'h3c0e: x = 16'h b6a; 14'h3c0f: x = 16'h b68; 14'h3c10: x = 16'h b67; 14'h3c11: x = 16'h b65; 14'h3c12: x = 16'h b64; 14'h3c13: x = 16'h b62; 14'h3c14: x = 16'h b61; 14'h3c15: x = 16'h b5f; 14'h3c16: x = 16'h b5e; 14'h3c17: x = 16'h b5c; 14'h3c18: x = 16'h b5b; 14'h3c19: x = 16'h b59; 14'h3c1a: x = 16'h b58; 14'h3c1b: x = 16'h b56; 14'h3c1c: x = 16'h b55; 14'h3c1d: x = 16'h b53; 14'h3c1e: x = 16'h b52; 14'h3c1f: x = 16'h b50; 14'h3c20: x = 16'h b4f; 14'h3c21: x = 16'h b4d; 14'h3c22: x = 16'h b4c; 14'h3c23: x = 16'h b4a; 14'h3c24: x = 16'h b49; 14'h3c25: x = 16'h b47; 14'h3c26: x = 16'h b46; 14'h3c27: x = 16'h b44; 14'h3c28: x = 16'h b43; 14'h3c29: x = 16'h b41; 14'h3c2a: x = 16'h b40; 14'h3c2b: x = 16'h b3e; 14'h3c2c: x = 16'h b3d; 14'h3c2d: x = 16'h b3b; 14'h3c2e: x = 16'h b3a; 14'h3c2f: x = 16'h b38; 14'h3c30: x = 16'h b37; 14'h3c31: x = 16'h b35; 14'h3c32: x = 16'h b34; 14'h3c33: x = 16'h b32; 14'h3c34: x = 16'h b31; 14'h3c35: x = 16'h b2f; 14'h3c36: x = 16'h b2e; 14'h3c37: x = 16'h b2c; 14'h3c38: x = 16'h b2a; 14'h3c39: x = 16'h b29; 14'h3c3a: x = 16'h b27; 14'h3c3b: x = 16'h b26; 14'h3c3c: x = 16'h b24; 14'h3c3d: x = 16'h b23; 14'h3c3e: x = 16'h b21; 14'h3c3f: x = 16'h b20; 14'h3c40: x = 16'h b1e; 14'h3c41: x = 16'h b1d; 14'h3c42: x = 16'h b1b; 14'h3c43: x = 16'h b1a; 14'h3c44: x = 16'h b18; 14'h3c45: x = 16'h b17; 14'h3c46: x = 16'h b15; 14'h3c47: x = 16'h b14; 14'h3c48: x = 16'h b12; 14'h3c49: x = 16'h b10; 14'h3c4a: x = 16'h b0f; 14'h3c4b: x = 16'h b0d; 14'h3c4c: x = 16'h b0c; 14'h3c4d: x = 16'h b0a; 14'h3c4e: x = 16'h b09; 14'h3c4f: x = 16'h b07; 14'h3c50: x = 16'h b06; 14'h3c51: x = 16'h b04; 14'h3c52: x = 16'h b03; 14'h3c53: x = 16'h b01; 14'h3c54: x = 16'h b00; 14'h3c55: x = 16'h afe; 14'h3c56: x = 16'h afc; 14'h3c57: x = 16'h afb; 14'h3c58: x = 16'h af9; 14'h3c59: x = 16'h af8; 14'h3c5a: x = 16'h af6; 14'h3c5b: x = 16'h af5; 14'h3c5c: x = 16'h af3; 14'h3c5d: x = 16'h af2; 14'h3c5e: x = 16'h af0; 14'h3c5f: x = 16'h aef; 14'h3c60: x = 16'h aed; 14'h3c61: x = 16'h aeb; 14'h3c62: x = 16'h aea; 14'h3c63: x = 16'h ae8; 14'h3c64: x = 16'h ae7; 14'h3c65: x = 16'h ae5; 14'h3c66: x = 16'h ae4; 14'h3c67: x = 16'h ae2; 14'h3c68: x = 16'h ae1; 14'h3c69: x = 16'h adf; 14'h3c6a: x = 16'h add; 14'h3c6b: x = 16'h adc; 14'h3c6c: x = 16'h ada; 14'h3c6d: x = 16'h ad9; 14'h3c6e: x = 16'h ad7; 14'h3c6f: x = 16'h ad6; 14'h3c70: x = 16'h ad4; 14'h3c71: x = 16'h ad2; 14'h3c72: x = 16'h ad1; 14'h3c73: x = 16'h acf; 14'h3c74: x = 16'h ace; 14'h3c75: x = 16'h acc; 14'h3c76: x = 16'h acb; 14'h3c77: x = 16'h ac9; 14'h3c78: x = 16'h ac8; 14'h3c79: x = 16'h ac6; 14'h3c7a: x = 16'h ac4; 14'h3c7b: x = 16'h ac3; 14'h3c7c: x = 16'h ac1; 14'h3c7d: x = 16'h ac0; 14'h3c7e: x = 16'h abe; 14'h3c7f: x = 16'h abd; 14'h3c80: x = 16'h abb; 14'h3c81: x = 16'h ab9; 14'h3c82: x = 16'h ab8; 14'h3c83: x = 16'h ab6; 14'h3c84: x = 16'h ab5; 14'h3c85: x = 16'h ab3; 14'h3c86: x = 16'h ab1; 14'h3c87: x = 16'h ab0; 14'h3c88: x = 16'h aae; 14'h3c89: x = 16'h aad; 14'h3c8a: x = 16'h aab; 14'h3c8b: x = 16'h aaa; 14'h3c8c: x = 16'h aa8; 14'h3c8d: x = 16'h aa6; 14'h3c8e: x = 16'h aa5; 14'h3c8f: x = 16'h aa3; 14'h3c90: x = 16'h aa2; 14'h3c91: x = 16'h aa0; 14'h3c92: x = 16'h a9e; 14'h3c93: x = 16'h a9d; 14'h3c94: x = 16'h a9b; 14'h3c95: x = 16'h a9a; 14'h3c96: x = 16'h a98; 14'h3c97: x = 16'h a96; 14'h3c98: x = 16'h a95; 14'h3c99: x = 16'h a93; 14'h3c9a: x = 16'h a92; 14'h3c9b: x = 16'h a90; 14'h3c9c: x = 16'h a8e; 14'h3c9d: x = 16'h a8d; 14'h3c9e: x = 16'h a8b; 14'h3c9f: x = 16'h a8a; 14'h3ca0: x = 16'h a88; 14'h3ca1: x = 16'h a86; 14'h3ca2: x = 16'h a85; 14'h3ca3: x = 16'h a83; 14'h3ca4: x = 16'h a82; 14'h3ca5: x = 16'h a80; 14'h3ca6: x = 16'h a7e; 14'h3ca7: x = 16'h a7d; 14'h3ca8: x = 16'h a7b; 14'h3ca9: x = 16'h a7a; 14'h3caa: x = 16'h a78; 14'h3cab: x = 16'h a76; 14'h3cac: x = 16'h a75; 14'h3cad: x = 16'h a73; 14'h3cae: x = 16'h a72; 14'h3caf: x = 16'h a70; 14'h3cb0: x = 16'h a6e; 14'h3cb1: x = 16'h a6d; 14'h3cb2: x = 16'h a6b; 14'h3cb3: x = 16'h a69; 14'h3cb4: x = 16'h a68; 14'h3cb5: x = 16'h a66; 14'h3cb6: x = 16'h a65; 14'h3cb7: x = 16'h a63; 14'h3cb8: x = 16'h a61; 14'h3cb9: x = 16'h a60; 14'h3cba: x = 16'h a5e; 14'h3cbb: x = 16'h a5c; 14'h3cbc: x = 16'h a5b; 14'h3cbd: x = 16'h a59; 14'h3cbe: x = 16'h a58; 14'h3cbf: x = 16'h a56; 14'h3cc0: x = 16'h a54; 14'h3cc1: x = 16'h a53; 14'h3cc2: x = 16'h a51; 14'h3cc3: x = 16'h a4f; 14'h3cc4: x = 16'h a4e; 14'h3cc5: x = 16'h a4c; 14'h3cc6: x = 16'h a4a; 14'h3cc7: x = 16'h a49; 14'h3cc8: x = 16'h a47; 14'h3cc9: x = 16'h a46; 14'h3cca: x = 16'h a44; 14'h3ccb: x = 16'h a42; 14'h3ccc: x = 16'h a41; 14'h3ccd: x = 16'h a3f; 14'h3cce: x = 16'h a3d; 14'h3ccf: x = 16'h a3c; 14'h3cd0: x = 16'h a3a; 14'h3cd1: x = 16'h a38; 14'h3cd2: x = 16'h a37; 14'h3cd3: x = 16'h a35; 14'h3cd4: x = 16'h a33; 14'h3cd5: x = 16'h a32; 14'h3cd6: x = 16'h a30; 14'h3cd7: x = 16'h a2f; 14'h3cd8: x = 16'h a2d; 14'h3cd9: x = 16'h a2b; 14'h3cda: x = 16'h a2a; 14'h3cdb: x = 16'h a28; 14'h3cdc: x = 16'h a26; 14'h3cdd: x = 16'h a25; 14'h3cde: x = 16'h a23; 14'h3cdf: x = 16'h a21; 14'h3ce0: x = 16'h a20; 14'h3ce1: x = 16'h a1e; 14'h3ce2: x = 16'h a1c; 14'h3ce3: x = 16'h a1b; 14'h3ce4: x = 16'h a19; 14'h3ce5: x = 16'h a17; 14'h3ce6: x = 16'h a16; 14'h3ce7: x = 16'h a14; 14'h3ce8: x = 16'h a12; 14'h3ce9: x = 16'h a11; 14'h3cea: x = 16'h a0f; 14'h3ceb: x = 16'h a0d; 14'h3cec: x = 16'h a0c; 14'h3ced: x = 16'h a0a; 14'h3cee: x = 16'h a08; 14'h3cef: x = 16'h a07; 14'h3cf0: x = 16'h a05; 14'h3cf1: x = 16'h a03; 14'h3cf2: x = 16'h a02; 14'h3cf3: x = 16'h a00; 14'h3cf4: x = 16'h 9fe; 14'h3cf5: x = 16'h 9fd; 14'h3cf6: x = 16'h 9fb; 14'h3cf7: x = 16'h 9f9; 14'h3cf8: x = 16'h 9f7; 14'h3cf9: x = 16'h 9f6; 14'h3cfa: x = 16'h 9f4; 14'h3cfb: x = 16'h 9f2; 14'h3cfc: x = 16'h 9f1; 14'h3cfd: x = 16'h 9ef; 14'h3cfe: x = 16'h 9ed; 14'h3cff: x = 16'h 9ec; 14'h3d00: x = 16'h 9ea; 14'h3d01: x = 16'h 9e8; 14'h3d02: x = 16'h 9e7; 14'h3d03: x = 16'h 9e5; 14'h3d04: x = 16'h 9e3; 14'h3d05: x = 16'h 9e1; 14'h3d06: x = 16'h 9e0; 14'h3d07: x = 16'h 9de; 14'h3d08: x = 16'h 9dc; 14'h3d09: x = 16'h 9db; 14'h3d0a: x = 16'h 9d9; 14'h3d0b: x = 16'h 9d7; 14'h3d0c: x = 16'h 9d6; 14'h3d0d: x = 16'h 9d4; 14'h3d0e: x = 16'h 9d2; 14'h3d0f: x = 16'h 9d0; 14'h3d10: x = 16'h 9cf; 14'h3d11: x = 16'h 9cd; 14'h3d12: x = 16'h 9cb; 14'h3d13: x = 16'h 9ca; 14'h3d14: x = 16'h 9c8; 14'h3d15: x = 16'h 9c6; 14'h3d16: x = 16'h 9c4; 14'h3d17: x = 16'h 9c3; 14'h3d18: x = 16'h 9c1; 14'h3d19: x = 16'h 9bf; 14'h3d1a: x = 16'h 9be; 14'h3d1b: x = 16'h 9bc; 14'h3d1c: x = 16'h 9ba; 14'h3d1d: x = 16'h 9b8; 14'h3d1e: x = 16'h 9b7; 14'h3d1f: x = 16'h 9b5; 14'h3d20: x = 16'h 9b3; 14'h3d21: x = 16'h 9b2; 14'h3d22: x = 16'h 9b0; 14'h3d23: x = 16'h 9ae; 14'h3d24: x = 16'h 9ac; 14'h3d25: x = 16'h 9ab; 14'h3d26: x = 16'h 9a9; 14'h3d27: x = 16'h 9a7; 14'h3d28: x = 16'h 9a5; 14'h3d29: x = 16'h 9a4; 14'h3d2a: x = 16'h 9a2; 14'h3d2b: x = 16'h 9a0; 14'h3d2c: x = 16'h 99e; 14'h3d2d: x = 16'h 99d; 14'h3d2e: x = 16'h 99b; 14'h3d2f: x = 16'h 999; 14'h3d30: x = 16'h 997; 14'h3d31: x = 16'h 996; 14'h3d32: x = 16'h 994; 14'h3d33: x = 16'h 992; 14'h3d34: x = 16'h 990; 14'h3d35: x = 16'h 98f; 14'h3d36: x = 16'h 98d; 14'h3d37: x = 16'h 98b; 14'h3d38: x = 16'h 989; 14'h3d39: x = 16'h 988; 14'h3d3a: x = 16'h 986; 14'h3d3b: x = 16'h 984; 14'h3d3c: x = 16'h 982; 14'h3d3d: x = 16'h 981; 14'h3d3e: x = 16'h 97f; 14'h3d3f: x = 16'h 97d; 14'h3d40: x = 16'h 97b; 14'h3d41: x = 16'h 97a; 14'h3d42: x = 16'h 978; 14'h3d43: x = 16'h 976; 14'h3d44: x = 16'h 974; 14'h3d45: x = 16'h 973; 14'h3d46: x = 16'h 971; 14'h3d47: x = 16'h 96f; 14'h3d48: x = 16'h 96d; 14'h3d49: x = 16'h 96b; 14'h3d4a: x = 16'h 96a; 14'h3d4b: x = 16'h 968; 14'h3d4c: x = 16'h 966; 14'h3d4d: x = 16'h 964; 14'h3d4e: x = 16'h 963; 14'h3d4f: x = 16'h 961; 14'h3d50: x = 16'h 95f; 14'h3d51: x = 16'h 95d; 14'h3d52: x = 16'h 95b; 14'h3d53: x = 16'h 95a; 14'h3d54: x = 16'h 958; 14'h3d55: x = 16'h 956; 14'h3d56: x = 16'h 954; 14'h3d57: x = 16'h 953; 14'h3d58: x = 16'h 951; 14'h3d59: x = 16'h 94f; 14'h3d5a: x = 16'h 94d; 14'h3d5b: x = 16'h 94b; 14'h3d5c: x = 16'h 94a; 14'h3d5d: x = 16'h 948; 14'h3d5e: x = 16'h 946; 14'h3d5f: x = 16'h 944; 14'h3d60: x = 16'h 942; 14'h3d61: x = 16'h 941; 14'h3d62: x = 16'h 93f; 14'h3d63: x = 16'h 93d; 14'h3d64: x = 16'h 93b; 14'h3d65: x = 16'h 939; 14'h3d66: x = 16'h 938; 14'h3d67: x = 16'h 936; 14'h3d68: x = 16'h 934; 14'h3d69: x = 16'h 932; 14'h3d6a: x = 16'h 930; 14'h3d6b: x = 16'h 92e; 14'h3d6c: x = 16'h 92d; 14'h3d6d: x = 16'h 92b; 14'h3d6e: x = 16'h 929; 14'h3d6f: x = 16'h 927; 14'h3d70: x = 16'h 925; 14'h3d71: x = 16'h 924; 14'h3d72: x = 16'h 922; 14'h3d73: x = 16'h 920; 14'h3d74: x = 16'h 91e; 14'h3d75: x = 16'h 91c; 14'h3d76: x = 16'h 91a; 14'h3d77: x = 16'h 919; 14'h3d78: x = 16'h 917; 14'h3d79: x = 16'h 915; 14'h3d7a: x = 16'h 913; 14'h3d7b: x = 16'h 911; 14'h3d7c: x = 16'h 90f; 14'h3d7d: x = 16'h 90e; 14'h3d7e: x = 16'h 90c; 14'h3d7f: x = 16'h 90a; 14'h3d80: x = 16'h 908; 14'h3d81: x = 16'h 906; 14'h3d82: x = 16'h 904; 14'h3d83: x = 16'h 903; 14'h3d84: x = 16'h 901; 14'h3d85: x = 16'h 8ff; 14'h3d86: x = 16'h 8fd; 14'h3d87: x = 16'h 8fb; 14'h3d88: x = 16'h 8f9; 14'h3d89: x = 16'h 8f7; 14'h3d8a: x = 16'h 8f6; 14'h3d8b: x = 16'h 8f4; 14'h3d8c: x = 16'h 8f2; 14'h3d8d: x = 16'h 8f0; 14'h3d8e: x = 16'h 8ee; 14'h3d8f: x = 16'h 8ec; 14'h3d90: x = 16'h 8ea; 14'h3d91: x = 16'h 8e9; 14'h3d92: x = 16'h 8e7; 14'h3d93: x = 16'h 8e5; 14'h3d94: x = 16'h 8e3; 14'h3d95: x = 16'h 8e1; 14'h3d96: x = 16'h 8df; 14'h3d97: x = 16'h 8dd; 14'h3d98: x = 16'h 8db; 14'h3d99: x = 16'h 8da; 14'h3d9a: x = 16'h 8d8; 14'h3d9b: x = 16'h 8d6; 14'h3d9c: x = 16'h 8d4; 14'h3d9d: x = 16'h 8d2; 14'h3d9e: x = 16'h 8d0; 14'h3d9f: x = 16'h 8ce; 14'h3da0: x = 16'h 8cc; 14'h3da1: x = 16'h 8ca; 14'h3da2: x = 16'h 8c9; 14'h3da3: x = 16'h 8c7; 14'h3da4: x = 16'h 8c5; 14'h3da5: x = 16'h 8c3; 14'h3da6: x = 16'h 8c1; 14'h3da7: x = 16'h 8bf; 14'h3da8: x = 16'h 8bd; 14'h3da9: x = 16'h 8bb; 14'h3daa: x = 16'h 8b9; 14'h3dab: x = 16'h 8b8; 14'h3dac: x = 16'h 8b6; 14'h3dad: x = 16'h 8b4; 14'h3dae: x = 16'h 8b2; 14'h3daf: x = 16'h 8b0; 14'h3db0: x = 16'h 8ae; 14'h3db1: x = 16'h 8ac; 14'h3db2: x = 16'h 8aa; 14'h3db3: x = 16'h 8a8; 14'h3db4: x = 16'h 8a6; 14'h3db5: x = 16'h 8a4; 14'h3db6: x = 16'h 8a2; 14'h3db7: x = 16'h 8a1; 14'h3db8: x = 16'h 89f; 14'h3db9: x = 16'h 89d; 14'h3dba: x = 16'h 89b; 14'h3dbb: x = 16'h 899; 14'h3dbc: x = 16'h 897; 14'h3dbd: x = 16'h 895; 14'h3dbe: x = 16'h 893; 14'h3dbf: x = 16'h 891; 14'h3dc0: x = 16'h 88f; 14'h3dc1: x = 16'h 88d; 14'h3dc2: x = 16'h 88b; 14'h3dc3: x = 16'h 889; 14'h3dc4: x = 16'h 887; 14'h3dc5: x = 16'h 885; 14'h3dc6: x = 16'h 884; 14'h3dc7: x = 16'h 882; 14'h3dc8: x = 16'h 880; 14'h3dc9: x = 16'h 87e; 14'h3dca: x = 16'h 87c; 14'h3dcb: x = 16'h 87a; 14'h3dcc: x = 16'h 878; 14'h3dcd: x = 16'h 876; 14'h3dce: x = 16'h 874; 14'h3dcf: x = 16'h 872; 14'h3dd0: x = 16'h 870; 14'h3dd1: x = 16'h 86e; 14'h3dd2: x = 16'h 86c; 14'h3dd3: x = 16'h 86a; 14'h3dd4: x = 16'h 868; 14'h3dd5: x = 16'h 866; 14'h3dd6: x = 16'h 864; 14'h3dd7: x = 16'h 862; 14'h3dd8: x = 16'h 860; 14'h3dd9: x = 16'h 85e; 14'h3dda: x = 16'h 85c; 14'h3ddb: x = 16'h 85a; 14'h3ddc: x = 16'h 858; 14'h3ddd: x = 16'h 856; 14'h3dde: x = 16'h 854; 14'h3ddf: x = 16'h 852; 14'h3de0: x = 16'h 850; 14'h3de1: x = 16'h 84e; 14'h3de2: x = 16'h 84c; 14'h3de3: x = 16'h 84a; 14'h3de4: x = 16'h 848; 14'h3de5: x = 16'h 846; 14'h3de6: x = 16'h 844; 14'h3de7: x = 16'h 842; 14'h3de8: x = 16'h 840; 14'h3de9: x = 16'h 83e; 14'h3dea: x = 16'h 83c; 14'h3deb: x = 16'h 83a; 14'h3dec: x = 16'h 838; 14'h3ded: x = 16'h 836; 14'h3dee: x = 16'h 834; 14'h3def: x = 16'h 832; 14'h3df0: x = 16'h 830; 14'h3df1: x = 16'h 82e; 14'h3df2: x = 16'h 82c; 14'h3df3: x = 16'h 82a; 14'h3df4: x = 16'h 828; 14'h3df5: x = 16'h 826; 14'h3df6: x = 16'h 824; 14'h3df7: x = 16'h 822; 14'h3df8: x = 16'h 820; 14'h3df9: x = 16'h 81e; 14'h3dfa: x = 16'h 81c; 14'h3dfb: x = 16'h 81a; 14'h3dfc: x = 16'h 818; 14'h3dfd: x = 16'h 816; 14'h3dfe: x = 16'h 814; 14'h3dff: x = 16'h 812; 14'h3e00: x = 16'h 810; 14'h3e01: x = 16'h 80e; 14'h3e02: x = 16'h 80c; 14'h3e03: x = 16'h 80a; 14'h3e04: x = 16'h 808; 14'h3e05: x = 16'h 806; 14'h3e06: x = 16'h 803; 14'h3e07: x = 16'h 801; 14'h3e08: x = 16'h 7ff; 14'h3e09: x = 16'h 7fd; 14'h3e0a: x = 16'h 7fb; 14'h3e0b: x = 16'h 7f9; 14'h3e0c: x = 16'h 7f7; 14'h3e0d: x = 16'h 7f5; 14'h3e0e: x = 16'h 7f3; 14'h3e0f: x = 16'h 7f1; 14'h3e10: x = 16'h 7ef; 14'h3e11: x = 16'h 7ed; 14'h3e12: x = 16'h 7eb; 14'h3e13: x = 16'h 7e9; 14'h3e14: x = 16'h 7e6; 14'h3e15: x = 16'h 7e4; 14'h3e16: x = 16'h 7e2; 14'h3e17: x = 16'h 7e0; 14'h3e18: x = 16'h 7de; 14'h3e19: x = 16'h 7dc; 14'h3e1a: x = 16'h 7da; 14'h3e1b: x = 16'h 7d8; 14'h3e1c: x = 16'h 7d6; 14'h3e1d: x = 16'h 7d4; 14'h3e1e: x = 16'h 7d1; 14'h3e1f: x = 16'h 7cf; 14'h3e20: x = 16'h 7cd; 14'h3e21: x = 16'h 7cb; 14'h3e22: x = 16'h 7c9; 14'h3e23: x = 16'h 7c7; 14'h3e24: x = 16'h 7c5; 14'h3e25: x = 16'h 7c3; 14'h3e26: x = 16'h 7c1; 14'h3e27: x = 16'h 7be; 14'h3e28: x = 16'h 7bc; 14'h3e29: x = 16'h 7ba; 14'h3e2a: x = 16'h 7b8; 14'h3e2b: x = 16'h 7b6; 14'h3e2c: x = 16'h 7b4; 14'h3e2d: x = 16'h 7b2; 14'h3e2e: x = 16'h 7af; 14'h3e2f: x = 16'h 7ad; 14'h3e30: x = 16'h 7ab; 14'h3e31: x = 16'h 7a9; 14'h3e32: x = 16'h 7a7; 14'h3e33: x = 16'h 7a5; 14'h3e34: x = 16'h 7a3; 14'h3e35: x = 16'h 7a0; 14'h3e36: x = 16'h 79e; 14'h3e37: x = 16'h 79c; 14'h3e38: x = 16'h 79a; 14'h3e39: x = 16'h 798; 14'h3e3a: x = 16'h 796; 14'h3e3b: x = 16'h 793; 14'h3e3c: x = 16'h 791; 14'h3e3d: x = 16'h 78f; 14'h3e3e: x = 16'h 78d; 14'h3e3f: x = 16'h 78b; 14'h3e40: x = 16'h 789; 14'h3e41: x = 16'h 786; 14'h3e42: x = 16'h 784; 14'h3e43: x = 16'h 782; 14'h3e44: x = 16'h 780; 14'h3e45: x = 16'h 77e; 14'h3e46: x = 16'h 77b; 14'h3e47: x = 16'h 779; 14'h3e48: x = 16'h 777; 14'h3e49: x = 16'h 775; 14'h3e4a: x = 16'h 773; 14'h3e4b: x = 16'h 770; 14'h3e4c: x = 16'h 76e; 14'h3e4d: x = 16'h 76c; 14'h3e4e: x = 16'h 76a; 14'h3e4f: x = 16'h 768; 14'h3e50: x = 16'h 765; 14'h3e51: x = 16'h 763; 14'h3e52: x = 16'h 761; 14'h3e53: x = 16'h 75f; 14'h3e54: x = 16'h 75c; 14'h3e55: x = 16'h 75a; 14'h3e56: x = 16'h 758; 14'h3e57: x = 16'h 756; 14'h3e58: x = 16'h 753; 14'h3e59: x = 16'h 751; 14'h3e5a: x = 16'h 74f; 14'h3e5b: x = 16'h 74d; 14'h3e5c: x = 16'h 74a; 14'h3e5d: x = 16'h 748; 14'h3e5e: x = 16'h 746; 14'h3e5f: x = 16'h 744; 14'h3e60: x = 16'h 741; 14'h3e61: x = 16'h 73f; 14'h3e62: x = 16'h 73d; 14'h3e63: x = 16'h 73b; 14'h3e64: x = 16'h 738; 14'h3e65: x = 16'h 736; 14'h3e66: x = 16'h 734; 14'h3e67: x = 16'h 732; 14'h3e68: x = 16'h 72f; 14'h3e69: x = 16'h 72d; 14'h3e6a: x = 16'h 72b; 14'h3e6b: x = 16'h 728; 14'h3e6c: x = 16'h 726; 14'h3e6d: x = 16'h 724; 14'h3e6e: x = 16'h 721; 14'h3e6f: x = 16'h 71f; 14'h3e70: x = 16'h 71d; 14'h3e71: x = 16'h 71b; 14'h3e72: x = 16'h 718; 14'h3e73: x = 16'h 716; 14'h3e74: x = 16'h 714; 14'h3e75: x = 16'h 711; 14'h3e76: x = 16'h 70f; 14'h3e77: x = 16'h 70d; 14'h3e78: x = 16'h 70a; 14'h3e79: x = 16'h 708; 14'h3e7a: x = 16'h 706; 14'h3e7b: x = 16'h 703; 14'h3e7c: x = 16'h 701; 14'h3e7d: x = 16'h 6ff; 14'h3e7e: x = 16'h 6fc; 14'h3e7f: x = 16'h 6fa; 14'h3e80: x = 16'h 6f8; 14'h3e81: x = 16'h 6f5; 14'h3e82: x = 16'h 6f3; 14'h3e83: x = 16'h 6f1; 14'h3e84: x = 16'h 6ee; 14'h3e85: x = 16'h 6ec; 14'h3e86: x = 16'h 6e9; 14'h3e87: x = 16'h 6e7; 14'h3e88: x = 16'h 6e5; 14'h3e89: x = 16'h 6e2; 14'h3e8a: x = 16'h 6e0; 14'h3e8b: x = 16'h 6de; 14'h3e8c: x = 16'h 6db; 14'h3e8d: x = 16'h 6d9; 14'h3e8e: x = 16'h 6d6; 14'h3e8f: x = 16'h 6d4; 14'h3e90: x = 16'h 6d2; 14'h3e91: x = 16'h 6cf; 14'h3e92: x = 16'h 6cd; 14'h3e93: x = 16'h 6ca; 14'h3e94: x = 16'h 6c8; 14'h3e95: x = 16'h 6c6; 14'h3e96: x = 16'h 6c3; 14'h3e97: x = 16'h 6c1; 14'h3e98: x = 16'h 6be; 14'h3e99: x = 16'h 6bc; 14'h3e9a: x = 16'h 6b9; 14'h3e9b: x = 16'h 6b7; 14'h3e9c: x = 16'h 6b5; 14'h3e9d: x = 16'h 6b2; 14'h3e9e: x = 16'h 6b0; 14'h3e9f: x = 16'h 6ad; 14'h3ea0: x = 16'h 6ab; 14'h3ea1: x = 16'h 6a8; 14'h3ea2: x = 16'h 6a6; 14'h3ea3: x = 16'h 6a3; 14'h3ea4: x = 16'h 6a1; 14'h3ea5: x = 16'h 69f; 14'h3ea6: x = 16'h 69c; 14'h3ea7: x = 16'h 69a; 14'h3ea8: x = 16'h 697; 14'h3ea9: x = 16'h 695; 14'h3eaa: x = 16'h 692; 14'h3eab: x = 16'h 690; 14'h3eac: x = 16'h 68d; 14'h3ead: x = 16'h 68b; 14'h3eae: x = 16'h 688; 14'h3eaf: x = 16'h 686; 14'h3eb0: x = 16'h 683; 14'h3eb1: x = 16'h 681; 14'h3eb2: x = 16'h 67e; 14'h3eb3: x = 16'h 67c; 14'h3eb4: x = 16'h 679; 14'h3eb5: x = 16'h 677; 14'h3eb6: x = 16'h 674; 14'h3eb7: x = 16'h 672; 14'h3eb8: x = 16'h 66f; 14'h3eb9: x = 16'h 66c; 14'h3eba: x = 16'h 66a; 14'h3ebb: x = 16'h 667; 14'h3ebc: x = 16'h 665; 14'h3ebd: x = 16'h 662; 14'h3ebe: x = 16'h 660; 14'h3ebf: x = 16'h 65d; 14'h3ec0: x = 16'h 65b; 14'h3ec1: x = 16'h 658; 14'h3ec2: x = 16'h 655; 14'h3ec3: x = 16'h 653; 14'h3ec4: x = 16'h 650; 14'h3ec5: x = 16'h 64e; 14'h3ec6: x = 16'h 64b; 14'h3ec7: x = 16'h 649; 14'h3ec8: x = 16'h 646; 14'h3ec9: x = 16'h 643; 14'h3eca: x = 16'h 641; 14'h3ecb: x = 16'h 63e; 14'h3ecc: x = 16'h 63b; 14'h3ecd: x = 16'h 639; 14'h3ece: x = 16'h 636; 14'h3ecf: x = 16'h 634; 14'h3ed0: x = 16'h 631; 14'h3ed1: x = 16'h 62e; 14'h3ed2: x = 16'h 62c; 14'h3ed3: x = 16'h 629; 14'h3ed4: x = 16'h 626; 14'h3ed5: x = 16'h 624; 14'h3ed6: x = 16'h 621; 14'h3ed7: x = 16'h 61e; 14'h3ed8: x = 16'h 61c; 14'h3ed9: x = 16'h 619; 14'h3eda: x = 16'h 616; 14'h3edb: x = 16'h 614; 14'h3edc: x = 16'h 611; 14'h3edd: x = 16'h 60e; 14'h3ede: x = 16'h 60c; 14'h3edf: x = 16'h 609; 14'h3ee0: x = 16'h 606; 14'h3ee1: x = 16'h 604; 14'h3ee2: x = 16'h 601; 14'h3ee3: x = 16'h 5fe; 14'h3ee4: x = 16'h 5fb; 14'h3ee5: x = 16'h 5f9; 14'h3ee6: x = 16'h 5f6; 14'h3ee7: x = 16'h 5f3; 14'h3ee8: x = 16'h 5f1; 14'h3ee9: x = 16'h 5ee; 14'h3eea: x = 16'h 5eb; 14'h3eeb: x = 16'h 5e8; 14'h3eec: x = 16'h 5e6; 14'h3eed: x = 16'h 5e3; 14'h3eee: x = 16'h 5e0; 14'h3eef: x = 16'h 5dd; 14'h3ef0: x = 16'h 5da; 14'h3ef1: x = 16'h 5d8; 14'h3ef2: x = 16'h 5d5; 14'h3ef3: x = 16'h 5d2; 14'h3ef4: x = 16'h 5cf; 14'h3ef5: x = 16'h 5cd; 14'h3ef6: x = 16'h 5ca; 14'h3ef7: x = 16'h 5c7; 14'h3ef8: x = 16'h 5c4; 14'h3ef9: x = 16'h 5c1; 14'h3efa: x = 16'h 5be; 14'h3efb: x = 16'h 5bc; 14'h3efc: x = 16'h 5b9; 14'h3efd: x = 16'h 5b6; 14'h3efe: x = 16'h 5b3; 14'h3eff: x = 16'h 5b0; 14'h3f00: x = 16'h 5ad; 14'h3f01: x = 16'h 5aa; 14'h3f02: x = 16'h 5a8; 14'h3f03: x = 16'h 5a5; 14'h3f04: x = 16'h 5a2; 14'h3f05: x = 16'h 59f; 14'h3f06: x = 16'h 59c; 14'h3f07: x = 16'h 599; 14'h3f08: x = 16'h 596; 14'h3f09: x = 16'h 593; 14'h3f0a: x = 16'h 590; 14'h3f0b: x = 16'h 58e; 14'h3f0c: x = 16'h 58b; 14'h3f0d: x = 16'h 588; 14'h3f0e: x = 16'h 585; 14'h3f0f: x = 16'h 582; 14'h3f10: x = 16'h 57f; 14'h3f11: x = 16'h 57c; 14'h3f12: x = 16'h 579; 14'h3f13: x = 16'h 576; 14'h3f14: x = 16'h 573; 14'h3f15: x = 16'h 570; 14'h3f16: x = 16'h 56d; 14'h3f17: x = 16'h 56a; 14'h3f18: x = 16'h 567; 14'h3f19: x = 16'h 564; 14'h3f1a: x = 16'h 561; 14'h3f1b: x = 16'h 55e; 14'h3f1c: x = 16'h 55b; 14'h3f1d: x = 16'h 558; 14'h3f1e: x = 16'h 555; 14'h3f1f: x = 16'h 552; 14'h3f20: x = 16'h 54f; 14'h3f21: x = 16'h 54c; 14'h3f22: x = 16'h 549; 14'h3f23: x = 16'h 546; 14'h3f24: x = 16'h 543; 14'h3f25: x = 16'h 53f; 14'h3f26: x = 16'h 53c; 14'h3f27: x = 16'h 539; 14'h3f28: x = 16'h 536; 14'h3f29: x = 16'h 533; 14'h3f2a: x = 16'h 530; 14'h3f2b: x = 16'h 52d; 14'h3f2c: x = 16'h 52a; 14'h3f2d: x = 16'h 526; 14'h3f2e: x = 16'h 523; 14'h3f2f: x = 16'h 520; 14'h3f30: x = 16'h 51d; 14'h3f31: x = 16'h 51a; 14'h3f32: x = 16'h 517; 14'h3f33: x = 16'h 513; 14'h3f34: x = 16'h 510; 14'h3f35: x = 16'h 50d; 14'h3f36: x = 16'h 50a; 14'h3f37: x = 16'h 507; 14'h3f38: x = 16'h 503; 14'h3f39: x = 16'h 500; 14'h3f3a: x = 16'h 4fd; 14'h3f3b: x = 16'h 4fa; 14'h3f3c: x = 16'h 4f6; 14'h3f3d: x = 16'h 4f3; 14'h3f3e: x = 16'h 4f0; 14'h3f3f: x = 16'h 4ed; 14'h3f40: x = 16'h 4e9; 14'h3f41: x = 16'h 4e6; 14'h3f42: x = 16'h 4e3; 14'h3f43: x = 16'h 4df; 14'h3f44: x = 16'h 4dc; 14'h3f45: x = 16'h 4d9; 14'h3f46: x = 16'h 4d5; 14'h3f47: x = 16'h 4d2; 14'h3f48: x = 16'h 4cf; 14'h3f49: x = 16'h 4cb; 14'h3f4a: x = 16'h 4c8; 14'h3f4b: x = 16'h 4c5; 14'h3f4c: x = 16'h 4c1; 14'h3f4d: x = 16'h 4be; 14'h3f4e: x = 16'h 4ba; 14'h3f4f: x = 16'h 4b7; 14'h3f50: x = 16'h 4b3; 14'h3f51: x = 16'h 4b0; 14'h3f52: x = 16'h 4ad; 14'h3f53: x = 16'h 4a9; 14'h3f54: x = 16'h 4a6; 14'h3f55: x = 16'h 4a2; 14'h3f56: x = 16'h 49f; 14'h3f57: x = 16'h 49b; 14'h3f58: x = 16'h 498; 14'h3f59: x = 16'h 494; 14'h3f5a: x = 16'h 491; 14'h3f5b: x = 16'h 48d; 14'h3f5c: x = 16'h 48a; 14'h3f5d: x = 16'h 486; 14'h3f5e: x = 16'h 482; 14'h3f5f: x = 16'h 47f; 14'h3f60: x = 16'h 47b; 14'h3f61: x = 16'h 478; 14'h3f62: x = 16'h 474; 14'h3f63: x = 16'h 470; 14'h3f64: x = 16'h 46d; 14'h3f65: x = 16'h 469; 14'h3f66: x = 16'h 465; 14'h3f67: x = 16'h 462; 14'h3f68: x = 16'h 45e; 14'h3f69: x = 16'h 45a; 14'h3f6a: x = 16'h 457; 14'h3f6b: x = 16'h 453; 14'h3f6c: x = 16'h 44f; 14'h3f6d: x = 16'h 44b; 14'h3f6e: x = 16'h 448; 14'h3f6f: x = 16'h 444; 14'h3f70: x = 16'h 440; 14'h3f71: x = 16'h 43c; 14'h3f72: x = 16'h 438; 14'h3f73: x = 16'h 435; 14'h3f74: x = 16'h 431; 14'h3f75: x = 16'h 42d; 14'h3f76: x = 16'h 429; 14'h3f77: x = 16'h 425; 14'h3f78: x = 16'h 421; 14'h3f79: x = 16'h 41d; 14'h3f7a: x = 16'h 419; 14'h3f7b: x = 16'h 415; 14'h3f7c: x = 16'h 411; 14'h3f7d: x = 16'h 40e; 14'h3f7e: x = 16'h 40a; 14'h3f7f: x = 16'h 406; 14'h3f80: x = 16'h 402; 14'h3f81: x = 16'h 3fd; 14'h3f82: x = 16'h 3f9; 14'h3f83: x = 16'h 3f5; 14'h3f84: x = 16'h 3f1; 14'h3f85: x = 16'h 3ed; 14'h3f86: x = 16'h 3e9; 14'h3f87: x = 16'h 3e5; 14'h3f88: x = 16'h 3e1; 14'h3f89: x = 16'h 3dd; 14'h3f8a: x = 16'h 3d8; 14'h3f8b: x = 16'h 3d4; 14'h3f8c: x = 16'h 3d0; 14'h3f8d: x = 16'h 3cc; 14'h3f8e: x = 16'h 3c8; 14'h3f8f: x = 16'h 3c3; 14'h3f90: x = 16'h 3bf; 14'h3f91: x = 16'h 3bb; 14'h3f92: x = 16'h 3b6; 14'h3f93: x = 16'h 3b2; 14'h3f94: x = 16'h 3ae; 14'h3f95: x = 16'h 3a9; 14'h3f96: x = 16'h 3a5; 14'h3f97: x = 16'h 3a0; 14'h3f98: x = 16'h 39c; 14'h3f99: x = 16'h 398; 14'h3f9a: x = 16'h 393; 14'h3f9b: x = 16'h 38f; 14'h3f9c: x = 16'h 38a; 14'h3f9d: x = 16'h 385; 14'h3f9e: x = 16'h 381; 14'h3f9f: x = 16'h 37c; 14'h3fa0: x = 16'h 378; 14'h3fa1: x = 16'h 373; 14'h3fa2: x = 16'h 36e; 14'h3fa3: x = 16'h 36a; 14'h3fa4: x = 16'h 365; 14'h3fa5: x = 16'h 360; 14'h3fa6: x = 16'h 35b; 14'h3fa7: x = 16'h 357; 14'h3fa8: x = 16'h 352; 14'h3fa9: x = 16'h 34d; 14'h3faa: x = 16'h 348; 14'h3fab: x = 16'h 343; 14'h3fac: x = 16'h 33e; 14'h3fad: x = 16'h 339; 14'h3fae: x = 16'h 334; 14'h3faf: x = 16'h 32f; 14'h3fb0: x = 16'h 32a; 14'h3fb1: x = 16'h 325; 14'h3fb2: x = 16'h 320; 14'h3fb3: x = 16'h 31b; 14'h3fb4: x = 16'h 315; 14'h3fb5: x = 16'h 310; 14'h3fb6: x = 16'h 30b; 14'h3fb7: x = 16'h 306; 14'h3fb8: x = 16'h 300; 14'h3fb9: x = 16'h 2fb; 14'h3fba: x = 16'h 2f6; 14'h3fbb: x = 16'h 2f0; 14'h3fbc: x = 16'h 2eb; 14'h3fbd: x = 16'h 2e5; 14'h3fbe: x = 16'h 2e0; 14'h3fbf: x = 16'h 2da; 14'h3fc0: x = 16'h 2d4; 14'h3fc1: x = 16'h 2cf; 14'h3fc2: x = 16'h 2c9; 14'h3fc3: x = 16'h 2c3; 14'h3fc4: x = 16'h 2bd; 14'h3fc5: x = 16'h 2b7; 14'h3fc6: x = 16'h 2b1; 14'h3fc7: x = 16'h 2ab; 14'h3fc8: x = 16'h 2a5; 14'h3fc9: x = 16'h 29f; 14'h3fca: x = 16'h 299; 14'h3fcb: x = 16'h 293; 14'h3fcc: x = 16'h 28d; 14'h3fcd: x = 16'h 286; 14'h3fce: x = 16'h 280; 14'h3fcf: x = 16'h 27a; 14'h3fd0: x = 16'h 273; 14'h3fd1: x = 16'h 26c; 14'h3fd2: x = 16'h 266; 14'h3fd3: x = 16'h 25f; 14'h3fd4: x = 16'h 258; 14'h3fd5: x = 16'h 251; 14'h3fd6: x = 16'h 24a; 14'h3fd7: x = 16'h 243; 14'h3fd8: x = 16'h 23c; 14'h3fd9: x = 16'h 235; 14'h3fda: x = 16'h 22e; 14'h3fdb: x = 16'h 226; 14'h3fdc: x = 16'h 21f; 14'h3fdd: x = 16'h 217; 14'h3fde: x = 16'h 210; 14'h3fdf: x = 16'h 208; 14'h3fe0: x = 16'h 200; 14'h3fe1: x = 16'h 1f8; 14'h3fe2: x = 16'h 1ef; 14'h3fe3: x = 16'h 1e7; 14'h3fe4: x = 16'h 1df; 14'h3fe5: x = 16'h 1d6; 14'h3fe6: x = 16'h 1cd; 14'h3fe7: x = 16'h 1c4; 14'h3fe8: x = 16'h 1bb; 14'h3fe9: x = 16'h 1b2; 14'h3fea: x = 16'h 1a8; 14'h3feb: x = 16'h 19e; 14'h3fec: x = 16'h 194; 14'h3fed: x = 16'h 18a; 14'h3fee: x = 16'h 180; 14'h3fef: x = 16'h 175; 14'h3ff0: x = 16'h 16a; 14'h3ff1: x = 16'h 15e; 14'h3ff2: x = 16'h 152; 14'h3ff3: x = 16'h 146; 14'h3ff4: x = 16'h 139; 14'h3ff5: x = 16'h 12c; 14'h3ff6: x = 16'h 11e; 14'h3ff7: x = 16'h 10f; 14'h3ff8: x = 16'h 100; 14'h3ff9: x = 16'h  ef; 14'h3ffa: x = 16'h  dd; 14'h3ffb: x = 16'h  ca; 14'h3ffc: x = 16'h  b5; 14'h3ffd: x = 16'h  9c; 14'h3ffe: x = 16'h  80; 14'h3fff: x = 16'h  5a; 
		default: x = 16'h0000;
		endcase
	end
endmodule

library ieee;
use ieee.std_logic_1164.all;

entity dot_disp1 is
port (
	clk : in std_logic;
	dot_data_00 : in std_logic_vector (6 downto 0);
	dot_data_01 : in std_logic_vector (6 downto 0);
	dot_data_02 : in std_logic_vector (6 downto 0);
	dot_data_03 : in std_logic_vector (6 downto 0);
	dot_data_04 : in std_logic_vector (6 downto 0);
	dot_data_05 : in std_logic_vector (6 downto 0);
	dot_data_06 : in std_logic_vector (6 downto 0);
	dot_data_07 : in std_logic_vector (6 downto 0);
	dot_data_08 : in std_logic_vector (6 downto 0);
	dot_data_09 : in std_logic_vector (6 downto 0);				
	dot_d : out std_logic_vector (6 downto 0);
	dot_scan : out std_logic_vector (9 downto 0);
	nreset  : in std_logic);
end dot_disp1;

architecture hb of dot_disp1 is
signal cnt_clk : integer range 0 to 9;
signal scan : std_logic_vector(9 downto 0);
begin

process(clk,nreset)
begin
	if nreset = '0' then
		cnt_clk <= 0;
	elsif clk'event and clk = '1' then
		if cnt_clk = 9 then
			cnt_clk <= 0;
		else
			cnt_clk <= cnt_clk + 1;
		end if;
	end if;
end process;

process(nreset,clk)
begin
	if nreset = '0' then
		scan <= "0000000001";
		dot_d <= "0000000";
	elsif clk'event and clk = '1' then
		if cnt_clk = 9 then
			scan <= "0000000001";
		else
			scan <= scan(8 downto 0) & '0';
		end if;
		
		case cnt_clk is
			when 0 =>
				dot_d <= dot_data_01;
			when 1 =>
				dot_d <= dot_data_02;
			when 2 =>
				dot_d <= dot_data_03;
			when 3 =>
				dot_d <= dot_data_04;
			when 4 =>
				dot_d <= dot_data_05;
			when 5 =>
				dot_d <= dot_data_06;
			when 6 =>
				dot_d <= dot_data_07;
			when 7 =>
				dot_d <= dot_data_08;
			when 8 =>
				dot_d <= dot_data_09;
			when 9 =>
				dot_d <= dot_data_00;
			when others => null;
		end case;
	end if;
end process;

	dot_scan <= scan;	

end hb;